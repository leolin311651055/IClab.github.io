# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : Img
#       Words            : 16384
#       Bits             : 8
#       Byte-Write       : 1
#       Aspect Ratio     : 8
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2025/05/22 14:41:46
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO Img
CLASS BLOCK ;
FOREIGN Img 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 1015.560 BY 764.400 ;
SYMMETRY x y r90 ;
SITE core_5040 ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 1014.440 752.980 1015.560 756.220 ;
  LAYER metal3 ;
  RECT 1014.440 752.980 1015.560 756.220 ;
  LAYER metal2 ;
  RECT 1014.440 752.980 1015.560 756.220 ;
  LAYER metal1 ;
  RECT 1014.440 752.980 1015.560 756.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 745.140 1015.560 748.380 ;
  LAYER metal3 ;
  RECT 1014.440 745.140 1015.560 748.380 ;
  LAYER metal2 ;
  RECT 1014.440 745.140 1015.560 748.380 ;
  LAYER metal1 ;
  RECT 1014.440 745.140 1015.560 748.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 737.300 1015.560 740.540 ;
  LAYER metal3 ;
  RECT 1014.440 737.300 1015.560 740.540 ;
  LAYER metal2 ;
  RECT 1014.440 737.300 1015.560 740.540 ;
  LAYER metal1 ;
  RECT 1014.440 737.300 1015.560 740.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 729.460 1015.560 732.700 ;
  LAYER metal3 ;
  RECT 1014.440 729.460 1015.560 732.700 ;
  LAYER metal2 ;
  RECT 1014.440 729.460 1015.560 732.700 ;
  LAYER metal1 ;
  RECT 1014.440 729.460 1015.560 732.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 721.620 1015.560 724.860 ;
  LAYER metal3 ;
  RECT 1014.440 721.620 1015.560 724.860 ;
  LAYER metal2 ;
  RECT 1014.440 721.620 1015.560 724.860 ;
  LAYER metal1 ;
  RECT 1014.440 721.620 1015.560 724.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 713.780 1015.560 717.020 ;
  LAYER metal3 ;
  RECT 1014.440 713.780 1015.560 717.020 ;
  LAYER metal2 ;
  RECT 1014.440 713.780 1015.560 717.020 ;
  LAYER metal1 ;
  RECT 1014.440 713.780 1015.560 717.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 674.580 1015.560 677.820 ;
  LAYER metal3 ;
  RECT 1014.440 674.580 1015.560 677.820 ;
  LAYER metal2 ;
  RECT 1014.440 674.580 1015.560 677.820 ;
  LAYER metal1 ;
  RECT 1014.440 674.580 1015.560 677.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 666.740 1015.560 669.980 ;
  LAYER metal3 ;
  RECT 1014.440 666.740 1015.560 669.980 ;
  LAYER metal2 ;
  RECT 1014.440 666.740 1015.560 669.980 ;
  LAYER metal1 ;
  RECT 1014.440 666.740 1015.560 669.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 658.900 1015.560 662.140 ;
  LAYER metal3 ;
  RECT 1014.440 658.900 1015.560 662.140 ;
  LAYER metal2 ;
  RECT 1014.440 658.900 1015.560 662.140 ;
  LAYER metal1 ;
  RECT 1014.440 658.900 1015.560 662.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 651.060 1015.560 654.300 ;
  LAYER metal3 ;
  RECT 1014.440 651.060 1015.560 654.300 ;
  LAYER metal2 ;
  RECT 1014.440 651.060 1015.560 654.300 ;
  LAYER metal1 ;
  RECT 1014.440 651.060 1015.560 654.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 643.220 1015.560 646.460 ;
  LAYER metal3 ;
  RECT 1014.440 643.220 1015.560 646.460 ;
  LAYER metal2 ;
  RECT 1014.440 643.220 1015.560 646.460 ;
  LAYER metal1 ;
  RECT 1014.440 643.220 1015.560 646.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 635.380 1015.560 638.620 ;
  LAYER metal3 ;
  RECT 1014.440 635.380 1015.560 638.620 ;
  LAYER metal2 ;
  RECT 1014.440 635.380 1015.560 638.620 ;
  LAYER metal1 ;
  RECT 1014.440 635.380 1015.560 638.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 596.180 1015.560 599.420 ;
  LAYER metal3 ;
  RECT 1014.440 596.180 1015.560 599.420 ;
  LAYER metal2 ;
  RECT 1014.440 596.180 1015.560 599.420 ;
  LAYER metal1 ;
  RECT 1014.440 596.180 1015.560 599.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 588.340 1015.560 591.580 ;
  LAYER metal3 ;
  RECT 1014.440 588.340 1015.560 591.580 ;
  LAYER metal2 ;
  RECT 1014.440 588.340 1015.560 591.580 ;
  LAYER metal1 ;
  RECT 1014.440 588.340 1015.560 591.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 580.500 1015.560 583.740 ;
  LAYER metal3 ;
  RECT 1014.440 580.500 1015.560 583.740 ;
  LAYER metal2 ;
  RECT 1014.440 580.500 1015.560 583.740 ;
  LAYER metal1 ;
  RECT 1014.440 580.500 1015.560 583.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 572.660 1015.560 575.900 ;
  LAYER metal3 ;
  RECT 1014.440 572.660 1015.560 575.900 ;
  LAYER metal2 ;
  RECT 1014.440 572.660 1015.560 575.900 ;
  LAYER metal1 ;
  RECT 1014.440 572.660 1015.560 575.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 564.820 1015.560 568.060 ;
  LAYER metal3 ;
  RECT 1014.440 564.820 1015.560 568.060 ;
  LAYER metal2 ;
  RECT 1014.440 564.820 1015.560 568.060 ;
  LAYER metal1 ;
  RECT 1014.440 564.820 1015.560 568.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 556.980 1015.560 560.220 ;
  LAYER metal3 ;
  RECT 1014.440 556.980 1015.560 560.220 ;
  LAYER metal2 ;
  RECT 1014.440 556.980 1015.560 560.220 ;
  LAYER metal1 ;
  RECT 1014.440 556.980 1015.560 560.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 517.780 1015.560 521.020 ;
  LAYER metal3 ;
  RECT 1014.440 517.780 1015.560 521.020 ;
  LAYER metal2 ;
  RECT 1014.440 517.780 1015.560 521.020 ;
  LAYER metal1 ;
  RECT 1014.440 517.780 1015.560 521.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 509.940 1015.560 513.180 ;
  LAYER metal3 ;
  RECT 1014.440 509.940 1015.560 513.180 ;
  LAYER metal2 ;
  RECT 1014.440 509.940 1015.560 513.180 ;
  LAYER metal1 ;
  RECT 1014.440 509.940 1015.560 513.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 502.100 1015.560 505.340 ;
  LAYER metal3 ;
  RECT 1014.440 502.100 1015.560 505.340 ;
  LAYER metal2 ;
  RECT 1014.440 502.100 1015.560 505.340 ;
  LAYER metal1 ;
  RECT 1014.440 502.100 1015.560 505.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 494.260 1015.560 497.500 ;
  LAYER metal3 ;
  RECT 1014.440 494.260 1015.560 497.500 ;
  LAYER metal2 ;
  RECT 1014.440 494.260 1015.560 497.500 ;
  LAYER metal1 ;
  RECT 1014.440 494.260 1015.560 497.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 486.420 1015.560 489.660 ;
  LAYER metal3 ;
  RECT 1014.440 486.420 1015.560 489.660 ;
  LAYER metal2 ;
  RECT 1014.440 486.420 1015.560 489.660 ;
  LAYER metal1 ;
  RECT 1014.440 486.420 1015.560 489.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 478.580 1015.560 481.820 ;
  LAYER metal3 ;
  RECT 1014.440 478.580 1015.560 481.820 ;
  LAYER metal2 ;
  RECT 1014.440 478.580 1015.560 481.820 ;
  LAYER metal1 ;
  RECT 1014.440 478.580 1015.560 481.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 439.380 1015.560 442.620 ;
  LAYER metal3 ;
  RECT 1014.440 439.380 1015.560 442.620 ;
  LAYER metal2 ;
  RECT 1014.440 439.380 1015.560 442.620 ;
  LAYER metal1 ;
  RECT 1014.440 439.380 1015.560 442.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 431.540 1015.560 434.780 ;
  LAYER metal3 ;
  RECT 1014.440 431.540 1015.560 434.780 ;
  LAYER metal2 ;
  RECT 1014.440 431.540 1015.560 434.780 ;
  LAYER metal1 ;
  RECT 1014.440 431.540 1015.560 434.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 423.700 1015.560 426.940 ;
  LAYER metal3 ;
  RECT 1014.440 423.700 1015.560 426.940 ;
  LAYER metal2 ;
  RECT 1014.440 423.700 1015.560 426.940 ;
  LAYER metal1 ;
  RECT 1014.440 423.700 1015.560 426.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 415.860 1015.560 419.100 ;
  LAYER metal3 ;
  RECT 1014.440 415.860 1015.560 419.100 ;
  LAYER metal2 ;
  RECT 1014.440 415.860 1015.560 419.100 ;
  LAYER metal1 ;
  RECT 1014.440 415.860 1015.560 419.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 408.020 1015.560 411.260 ;
  LAYER metal3 ;
  RECT 1014.440 408.020 1015.560 411.260 ;
  LAYER metal2 ;
  RECT 1014.440 408.020 1015.560 411.260 ;
  LAYER metal1 ;
  RECT 1014.440 408.020 1015.560 411.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 400.180 1015.560 403.420 ;
  LAYER metal3 ;
  RECT 1014.440 400.180 1015.560 403.420 ;
  LAYER metal2 ;
  RECT 1014.440 400.180 1015.560 403.420 ;
  LAYER metal1 ;
  RECT 1014.440 400.180 1015.560 403.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 360.980 1015.560 364.220 ;
  LAYER metal3 ;
  RECT 1014.440 360.980 1015.560 364.220 ;
  LAYER metal2 ;
  RECT 1014.440 360.980 1015.560 364.220 ;
  LAYER metal1 ;
  RECT 1014.440 360.980 1015.560 364.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 353.140 1015.560 356.380 ;
  LAYER metal3 ;
  RECT 1014.440 353.140 1015.560 356.380 ;
  LAYER metal2 ;
  RECT 1014.440 353.140 1015.560 356.380 ;
  LAYER metal1 ;
  RECT 1014.440 353.140 1015.560 356.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 345.300 1015.560 348.540 ;
  LAYER metal3 ;
  RECT 1014.440 345.300 1015.560 348.540 ;
  LAYER metal2 ;
  RECT 1014.440 345.300 1015.560 348.540 ;
  LAYER metal1 ;
  RECT 1014.440 345.300 1015.560 348.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 337.460 1015.560 340.700 ;
  LAYER metal3 ;
  RECT 1014.440 337.460 1015.560 340.700 ;
  LAYER metal2 ;
  RECT 1014.440 337.460 1015.560 340.700 ;
  LAYER metal1 ;
  RECT 1014.440 337.460 1015.560 340.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 329.620 1015.560 332.860 ;
  LAYER metal3 ;
  RECT 1014.440 329.620 1015.560 332.860 ;
  LAYER metal2 ;
  RECT 1014.440 329.620 1015.560 332.860 ;
  LAYER metal1 ;
  RECT 1014.440 329.620 1015.560 332.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 321.780 1015.560 325.020 ;
  LAYER metal3 ;
  RECT 1014.440 321.780 1015.560 325.020 ;
  LAYER metal2 ;
  RECT 1014.440 321.780 1015.560 325.020 ;
  LAYER metal1 ;
  RECT 1014.440 321.780 1015.560 325.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 282.580 1015.560 285.820 ;
  LAYER metal3 ;
  RECT 1014.440 282.580 1015.560 285.820 ;
  LAYER metal2 ;
  RECT 1014.440 282.580 1015.560 285.820 ;
  LAYER metal1 ;
  RECT 1014.440 282.580 1015.560 285.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 274.740 1015.560 277.980 ;
  LAYER metal3 ;
  RECT 1014.440 274.740 1015.560 277.980 ;
  LAYER metal2 ;
  RECT 1014.440 274.740 1015.560 277.980 ;
  LAYER metal1 ;
  RECT 1014.440 274.740 1015.560 277.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 266.900 1015.560 270.140 ;
  LAYER metal3 ;
  RECT 1014.440 266.900 1015.560 270.140 ;
  LAYER metal2 ;
  RECT 1014.440 266.900 1015.560 270.140 ;
  LAYER metal1 ;
  RECT 1014.440 266.900 1015.560 270.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 259.060 1015.560 262.300 ;
  LAYER metal3 ;
  RECT 1014.440 259.060 1015.560 262.300 ;
  LAYER metal2 ;
  RECT 1014.440 259.060 1015.560 262.300 ;
  LAYER metal1 ;
  RECT 1014.440 259.060 1015.560 262.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 251.220 1015.560 254.460 ;
  LAYER metal3 ;
  RECT 1014.440 251.220 1015.560 254.460 ;
  LAYER metal2 ;
  RECT 1014.440 251.220 1015.560 254.460 ;
  LAYER metal1 ;
  RECT 1014.440 251.220 1015.560 254.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 243.380 1015.560 246.620 ;
  LAYER metal3 ;
  RECT 1014.440 243.380 1015.560 246.620 ;
  LAYER metal2 ;
  RECT 1014.440 243.380 1015.560 246.620 ;
  LAYER metal1 ;
  RECT 1014.440 243.380 1015.560 246.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 204.180 1015.560 207.420 ;
  LAYER metal3 ;
  RECT 1014.440 204.180 1015.560 207.420 ;
  LAYER metal2 ;
  RECT 1014.440 204.180 1015.560 207.420 ;
  LAYER metal1 ;
  RECT 1014.440 204.180 1015.560 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 196.340 1015.560 199.580 ;
  LAYER metal3 ;
  RECT 1014.440 196.340 1015.560 199.580 ;
  LAYER metal2 ;
  RECT 1014.440 196.340 1015.560 199.580 ;
  LAYER metal1 ;
  RECT 1014.440 196.340 1015.560 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 188.500 1015.560 191.740 ;
  LAYER metal3 ;
  RECT 1014.440 188.500 1015.560 191.740 ;
  LAYER metal2 ;
  RECT 1014.440 188.500 1015.560 191.740 ;
  LAYER metal1 ;
  RECT 1014.440 188.500 1015.560 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 180.660 1015.560 183.900 ;
  LAYER metal3 ;
  RECT 1014.440 180.660 1015.560 183.900 ;
  LAYER metal2 ;
  RECT 1014.440 180.660 1015.560 183.900 ;
  LAYER metal1 ;
  RECT 1014.440 180.660 1015.560 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 172.820 1015.560 176.060 ;
  LAYER metal3 ;
  RECT 1014.440 172.820 1015.560 176.060 ;
  LAYER metal2 ;
  RECT 1014.440 172.820 1015.560 176.060 ;
  LAYER metal1 ;
  RECT 1014.440 172.820 1015.560 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 164.980 1015.560 168.220 ;
  LAYER metal3 ;
  RECT 1014.440 164.980 1015.560 168.220 ;
  LAYER metal2 ;
  RECT 1014.440 164.980 1015.560 168.220 ;
  LAYER metal1 ;
  RECT 1014.440 164.980 1015.560 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 125.780 1015.560 129.020 ;
  LAYER metal3 ;
  RECT 1014.440 125.780 1015.560 129.020 ;
  LAYER metal2 ;
  RECT 1014.440 125.780 1015.560 129.020 ;
  LAYER metal1 ;
  RECT 1014.440 125.780 1015.560 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 117.940 1015.560 121.180 ;
  LAYER metal3 ;
  RECT 1014.440 117.940 1015.560 121.180 ;
  LAYER metal2 ;
  RECT 1014.440 117.940 1015.560 121.180 ;
  LAYER metal1 ;
  RECT 1014.440 117.940 1015.560 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 110.100 1015.560 113.340 ;
  LAYER metal3 ;
  RECT 1014.440 110.100 1015.560 113.340 ;
  LAYER metal2 ;
  RECT 1014.440 110.100 1015.560 113.340 ;
  LAYER metal1 ;
  RECT 1014.440 110.100 1015.560 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 102.260 1015.560 105.500 ;
  LAYER metal3 ;
  RECT 1014.440 102.260 1015.560 105.500 ;
  LAYER metal2 ;
  RECT 1014.440 102.260 1015.560 105.500 ;
  LAYER metal1 ;
  RECT 1014.440 102.260 1015.560 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 94.420 1015.560 97.660 ;
  LAYER metal3 ;
  RECT 1014.440 94.420 1015.560 97.660 ;
  LAYER metal2 ;
  RECT 1014.440 94.420 1015.560 97.660 ;
  LAYER metal1 ;
  RECT 1014.440 94.420 1015.560 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 86.580 1015.560 89.820 ;
  LAYER metal3 ;
  RECT 1014.440 86.580 1015.560 89.820 ;
  LAYER metal2 ;
  RECT 1014.440 86.580 1015.560 89.820 ;
  LAYER metal1 ;
  RECT 1014.440 86.580 1015.560 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 47.380 1015.560 50.620 ;
  LAYER metal3 ;
  RECT 1014.440 47.380 1015.560 50.620 ;
  LAYER metal2 ;
  RECT 1014.440 47.380 1015.560 50.620 ;
  LAYER metal1 ;
  RECT 1014.440 47.380 1015.560 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 39.540 1015.560 42.780 ;
  LAYER metal3 ;
  RECT 1014.440 39.540 1015.560 42.780 ;
  LAYER metal2 ;
  RECT 1014.440 39.540 1015.560 42.780 ;
  LAYER metal1 ;
  RECT 1014.440 39.540 1015.560 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 31.700 1015.560 34.940 ;
  LAYER metal3 ;
  RECT 1014.440 31.700 1015.560 34.940 ;
  LAYER metal2 ;
  RECT 1014.440 31.700 1015.560 34.940 ;
  LAYER metal1 ;
  RECT 1014.440 31.700 1015.560 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 23.860 1015.560 27.100 ;
  LAYER metal3 ;
  RECT 1014.440 23.860 1015.560 27.100 ;
  LAYER metal2 ;
  RECT 1014.440 23.860 1015.560 27.100 ;
  LAYER metal1 ;
  RECT 1014.440 23.860 1015.560 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 16.020 1015.560 19.260 ;
  LAYER metal3 ;
  RECT 1014.440 16.020 1015.560 19.260 ;
  LAYER metal2 ;
  RECT 1014.440 16.020 1015.560 19.260 ;
  LAYER metal1 ;
  RECT 1014.440 16.020 1015.560 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 8.180 1015.560 11.420 ;
  LAYER metal3 ;
  RECT 1014.440 8.180 1015.560 11.420 ;
  LAYER metal2 ;
  RECT 1014.440 8.180 1015.560 11.420 ;
  LAYER metal1 ;
  RECT 1014.440 8.180 1015.560 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 752.980 1.120 756.220 ;
  LAYER metal3 ;
  RECT 0.000 752.980 1.120 756.220 ;
  LAYER metal2 ;
  RECT 0.000 752.980 1.120 756.220 ;
  LAYER metal1 ;
  RECT 0.000 752.980 1.120 756.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 745.140 1.120 748.380 ;
  LAYER metal3 ;
  RECT 0.000 745.140 1.120 748.380 ;
  LAYER metal2 ;
  RECT 0.000 745.140 1.120 748.380 ;
  LAYER metal1 ;
  RECT 0.000 745.140 1.120 748.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 737.300 1.120 740.540 ;
  LAYER metal3 ;
  RECT 0.000 737.300 1.120 740.540 ;
  LAYER metal2 ;
  RECT 0.000 737.300 1.120 740.540 ;
  LAYER metal1 ;
  RECT 0.000 737.300 1.120 740.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 729.460 1.120 732.700 ;
  LAYER metal3 ;
  RECT 0.000 729.460 1.120 732.700 ;
  LAYER metal2 ;
  RECT 0.000 729.460 1.120 732.700 ;
  LAYER metal1 ;
  RECT 0.000 729.460 1.120 732.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 721.620 1.120 724.860 ;
  LAYER metal3 ;
  RECT 0.000 721.620 1.120 724.860 ;
  LAYER metal2 ;
  RECT 0.000 721.620 1.120 724.860 ;
  LAYER metal1 ;
  RECT 0.000 721.620 1.120 724.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 713.780 1.120 717.020 ;
  LAYER metal3 ;
  RECT 0.000 713.780 1.120 717.020 ;
  LAYER metal2 ;
  RECT 0.000 713.780 1.120 717.020 ;
  LAYER metal1 ;
  RECT 0.000 713.780 1.120 717.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 674.580 1.120 677.820 ;
  LAYER metal3 ;
  RECT 0.000 674.580 1.120 677.820 ;
  LAYER metal2 ;
  RECT 0.000 674.580 1.120 677.820 ;
  LAYER metal1 ;
  RECT 0.000 674.580 1.120 677.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 666.740 1.120 669.980 ;
  LAYER metal3 ;
  RECT 0.000 666.740 1.120 669.980 ;
  LAYER metal2 ;
  RECT 0.000 666.740 1.120 669.980 ;
  LAYER metal1 ;
  RECT 0.000 666.740 1.120 669.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 658.900 1.120 662.140 ;
  LAYER metal3 ;
  RECT 0.000 658.900 1.120 662.140 ;
  LAYER metal2 ;
  RECT 0.000 658.900 1.120 662.140 ;
  LAYER metal1 ;
  RECT 0.000 658.900 1.120 662.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 651.060 1.120 654.300 ;
  LAYER metal3 ;
  RECT 0.000 651.060 1.120 654.300 ;
  LAYER metal2 ;
  RECT 0.000 651.060 1.120 654.300 ;
  LAYER metal1 ;
  RECT 0.000 651.060 1.120 654.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 643.220 1.120 646.460 ;
  LAYER metal3 ;
  RECT 0.000 643.220 1.120 646.460 ;
  LAYER metal2 ;
  RECT 0.000 643.220 1.120 646.460 ;
  LAYER metal1 ;
  RECT 0.000 643.220 1.120 646.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 635.380 1.120 638.620 ;
  LAYER metal3 ;
  RECT 0.000 635.380 1.120 638.620 ;
  LAYER metal2 ;
  RECT 0.000 635.380 1.120 638.620 ;
  LAYER metal1 ;
  RECT 0.000 635.380 1.120 638.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 596.180 1.120 599.420 ;
  LAYER metal3 ;
  RECT 0.000 596.180 1.120 599.420 ;
  LAYER metal2 ;
  RECT 0.000 596.180 1.120 599.420 ;
  LAYER metal1 ;
  RECT 0.000 596.180 1.120 599.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 588.340 1.120 591.580 ;
  LAYER metal3 ;
  RECT 0.000 588.340 1.120 591.580 ;
  LAYER metal2 ;
  RECT 0.000 588.340 1.120 591.580 ;
  LAYER metal1 ;
  RECT 0.000 588.340 1.120 591.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 580.500 1.120 583.740 ;
  LAYER metal3 ;
  RECT 0.000 580.500 1.120 583.740 ;
  LAYER metal2 ;
  RECT 0.000 580.500 1.120 583.740 ;
  LAYER metal1 ;
  RECT 0.000 580.500 1.120 583.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 572.660 1.120 575.900 ;
  LAYER metal3 ;
  RECT 0.000 572.660 1.120 575.900 ;
  LAYER metal2 ;
  RECT 0.000 572.660 1.120 575.900 ;
  LAYER metal1 ;
  RECT 0.000 572.660 1.120 575.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 564.820 1.120 568.060 ;
  LAYER metal3 ;
  RECT 0.000 564.820 1.120 568.060 ;
  LAYER metal2 ;
  RECT 0.000 564.820 1.120 568.060 ;
  LAYER metal1 ;
  RECT 0.000 564.820 1.120 568.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 556.980 1.120 560.220 ;
  LAYER metal3 ;
  RECT 0.000 556.980 1.120 560.220 ;
  LAYER metal2 ;
  RECT 0.000 556.980 1.120 560.220 ;
  LAYER metal1 ;
  RECT 0.000 556.980 1.120 560.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER metal3 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER metal2 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER metal1 ;
  RECT 0.000 517.780 1.120 521.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER metal3 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER metal2 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER metal1 ;
  RECT 0.000 509.940 1.120 513.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER metal3 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER metal2 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER metal1 ;
  RECT 0.000 502.100 1.120 505.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER metal3 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER metal2 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER metal1 ;
  RECT 0.000 494.260 1.120 497.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER metal3 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER metal2 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER metal1 ;
  RECT 0.000 486.420 1.120 489.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER metal3 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER metal2 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER metal1 ;
  RECT 0.000 478.580 1.120 481.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER metal3 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER metal2 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER metal1 ;
  RECT 0.000 439.380 1.120 442.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER metal3 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER metal2 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER metal1 ;
  RECT 0.000 431.540 1.120 434.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER metal3 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER metal2 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER metal1 ;
  RECT 0.000 423.700 1.120 426.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER metal3 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER metal2 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER metal1 ;
  RECT 0.000 415.860 1.120 419.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER metal3 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER metal2 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER metal1 ;
  RECT 0.000 408.020 1.120 411.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER metal3 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER metal2 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER metal1 ;
  RECT 0.000 400.180 1.120 403.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER metal3 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER metal2 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER metal1 ;
  RECT 0.000 360.980 1.120 364.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER metal3 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER metal2 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER metal1 ;
  RECT 0.000 353.140 1.120 356.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER metal3 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER metal2 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER metal1 ;
  RECT 0.000 345.300 1.120 348.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER metal3 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER metal2 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER metal1 ;
  RECT 0.000 337.460 1.120 340.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER metal3 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER metal2 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER metal1 ;
  RECT 0.000 329.620 1.120 332.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER metal3 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER metal2 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER metal1 ;
  RECT 0.000 321.780 1.120 325.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal3 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal2 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal1 ;
  RECT 0.000 282.580 1.120 285.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal3 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal2 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal1 ;
  RECT 0.000 274.740 1.120 277.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal3 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal2 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal1 ;
  RECT 0.000 266.900 1.120 270.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal3 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal2 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal1 ;
  RECT 0.000 259.060 1.120 262.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal3 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal2 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal1 ;
  RECT 0.000 251.220 1.120 254.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal3 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal2 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal1 ;
  RECT 0.000 243.380 1.120 246.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 997.360 763.280 1000.900 764.400 ;
  LAYER metal3 ;
  RECT 997.360 763.280 1000.900 764.400 ;
  LAYER metal2 ;
  RECT 997.360 763.280 1000.900 764.400 ;
  LAYER metal1 ;
  RECT 997.360 763.280 1000.900 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 988.680 763.280 992.220 764.400 ;
  LAYER metal3 ;
  RECT 988.680 763.280 992.220 764.400 ;
  LAYER metal2 ;
  RECT 988.680 763.280 992.220 764.400 ;
  LAYER metal1 ;
  RECT 988.680 763.280 992.220 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 980.000 763.280 983.540 764.400 ;
  LAYER metal3 ;
  RECT 980.000 763.280 983.540 764.400 ;
  LAYER metal2 ;
  RECT 980.000 763.280 983.540 764.400 ;
  LAYER metal1 ;
  RECT 980.000 763.280 983.540 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 971.320 763.280 974.860 764.400 ;
  LAYER metal3 ;
  RECT 971.320 763.280 974.860 764.400 ;
  LAYER metal2 ;
  RECT 971.320 763.280 974.860 764.400 ;
  LAYER metal1 ;
  RECT 971.320 763.280 974.860 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 962.640 763.280 966.180 764.400 ;
  LAYER metal3 ;
  RECT 962.640 763.280 966.180 764.400 ;
  LAYER metal2 ;
  RECT 962.640 763.280 966.180 764.400 ;
  LAYER metal1 ;
  RECT 962.640 763.280 966.180 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 919.240 763.280 922.780 764.400 ;
  LAYER metal3 ;
  RECT 919.240 763.280 922.780 764.400 ;
  LAYER metal2 ;
  RECT 919.240 763.280 922.780 764.400 ;
  LAYER metal1 ;
  RECT 919.240 763.280 922.780 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 910.560 763.280 914.100 764.400 ;
  LAYER metal3 ;
  RECT 910.560 763.280 914.100 764.400 ;
  LAYER metal2 ;
  RECT 910.560 763.280 914.100 764.400 ;
  LAYER metal1 ;
  RECT 910.560 763.280 914.100 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 901.880 763.280 905.420 764.400 ;
  LAYER metal3 ;
  RECT 901.880 763.280 905.420 764.400 ;
  LAYER metal2 ;
  RECT 901.880 763.280 905.420 764.400 ;
  LAYER metal1 ;
  RECT 901.880 763.280 905.420 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 893.200 763.280 896.740 764.400 ;
  LAYER metal3 ;
  RECT 893.200 763.280 896.740 764.400 ;
  LAYER metal2 ;
  RECT 893.200 763.280 896.740 764.400 ;
  LAYER metal1 ;
  RECT 893.200 763.280 896.740 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 884.520 763.280 888.060 764.400 ;
  LAYER metal3 ;
  RECT 884.520 763.280 888.060 764.400 ;
  LAYER metal2 ;
  RECT 884.520 763.280 888.060 764.400 ;
  LAYER metal1 ;
  RECT 884.520 763.280 888.060 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 875.840 763.280 879.380 764.400 ;
  LAYER metal3 ;
  RECT 875.840 763.280 879.380 764.400 ;
  LAYER metal2 ;
  RECT 875.840 763.280 879.380 764.400 ;
  LAYER metal1 ;
  RECT 875.840 763.280 879.380 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 832.440 763.280 835.980 764.400 ;
  LAYER metal3 ;
  RECT 832.440 763.280 835.980 764.400 ;
  LAYER metal2 ;
  RECT 832.440 763.280 835.980 764.400 ;
  LAYER metal1 ;
  RECT 832.440 763.280 835.980 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 823.760 763.280 827.300 764.400 ;
  LAYER metal3 ;
  RECT 823.760 763.280 827.300 764.400 ;
  LAYER metal2 ;
  RECT 823.760 763.280 827.300 764.400 ;
  LAYER metal1 ;
  RECT 823.760 763.280 827.300 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 815.080 763.280 818.620 764.400 ;
  LAYER metal3 ;
  RECT 815.080 763.280 818.620 764.400 ;
  LAYER metal2 ;
  RECT 815.080 763.280 818.620 764.400 ;
  LAYER metal1 ;
  RECT 815.080 763.280 818.620 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 806.400 763.280 809.940 764.400 ;
  LAYER metal3 ;
  RECT 806.400 763.280 809.940 764.400 ;
  LAYER metal2 ;
  RECT 806.400 763.280 809.940 764.400 ;
  LAYER metal1 ;
  RECT 806.400 763.280 809.940 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 797.720 763.280 801.260 764.400 ;
  LAYER metal3 ;
  RECT 797.720 763.280 801.260 764.400 ;
  LAYER metal2 ;
  RECT 797.720 763.280 801.260 764.400 ;
  LAYER metal1 ;
  RECT 797.720 763.280 801.260 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 789.040 763.280 792.580 764.400 ;
  LAYER metal3 ;
  RECT 789.040 763.280 792.580 764.400 ;
  LAYER metal2 ;
  RECT 789.040 763.280 792.580 764.400 ;
  LAYER metal1 ;
  RECT 789.040 763.280 792.580 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 745.640 763.280 749.180 764.400 ;
  LAYER metal3 ;
  RECT 745.640 763.280 749.180 764.400 ;
  LAYER metal2 ;
  RECT 745.640 763.280 749.180 764.400 ;
  LAYER metal1 ;
  RECT 745.640 763.280 749.180 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 736.960 763.280 740.500 764.400 ;
  LAYER metal3 ;
  RECT 736.960 763.280 740.500 764.400 ;
  LAYER metal2 ;
  RECT 736.960 763.280 740.500 764.400 ;
  LAYER metal1 ;
  RECT 736.960 763.280 740.500 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 728.280 763.280 731.820 764.400 ;
  LAYER metal3 ;
  RECT 728.280 763.280 731.820 764.400 ;
  LAYER metal2 ;
  RECT 728.280 763.280 731.820 764.400 ;
  LAYER metal1 ;
  RECT 728.280 763.280 731.820 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 719.600 763.280 723.140 764.400 ;
  LAYER metal3 ;
  RECT 719.600 763.280 723.140 764.400 ;
  LAYER metal2 ;
  RECT 719.600 763.280 723.140 764.400 ;
  LAYER metal1 ;
  RECT 719.600 763.280 723.140 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 710.920 763.280 714.460 764.400 ;
  LAYER metal3 ;
  RECT 710.920 763.280 714.460 764.400 ;
  LAYER metal2 ;
  RECT 710.920 763.280 714.460 764.400 ;
  LAYER metal1 ;
  RECT 710.920 763.280 714.460 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 702.240 763.280 705.780 764.400 ;
  LAYER metal3 ;
  RECT 702.240 763.280 705.780 764.400 ;
  LAYER metal2 ;
  RECT 702.240 763.280 705.780 764.400 ;
  LAYER metal1 ;
  RECT 702.240 763.280 705.780 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 658.840 763.280 662.380 764.400 ;
  LAYER metal3 ;
  RECT 658.840 763.280 662.380 764.400 ;
  LAYER metal2 ;
  RECT 658.840 763.280 662.380 764.400 ;
  LAYER metal1 ;
  RECT 658.840 763.280 662.380 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 650.160 763.280 653.700 764.400 ;
  LAYER metal3 ;
  RECT 650.160 763.280 653.700 764.400 ;
  LAYER metal2 ;
  RECT 650.160 763.280 653.700 764.400 ;
  LAYER metal1 ;
  RECT 650.160 763.280 653.700 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 641.480 763.280 645.020 764.400 ;
  LAYER metal3 ;
  RECT 641.480 763.280 645.020 764.400 ;
  LAYER metal2 ;
  RECT 641.480 763.280 645.020 764.400 ;
  LAYER metal1 ;
  RECT 641.480 763.280 645.020 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 632.800 763.280 636.340 764.400 ;
  LAYER metal3 ;
  RECT 632.800 763.280 636.340 764.400 ;
  LAYER metal2 ;
  RECT 632.800 763.280 636.340 764.400 ;
  LAYER metal1 ;
  RECT 632.800 763.280 636.340 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 624.120 763.280 627.660 764.400 ;
  LAYER metal3 ;
  RECT 624.120 763.280 627.660 764.400 ;
  LAYER metal2 ;
  RECT 624.120 763.280 627.660 764.400 ;
  LAYER metal1 ;
  RECT 624.120 763.280 627.660 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 615.440 763.280 618.980 764.400 ;
  LAYER metal3 ;
  RECT 615.440 763.280 618.980 764.400 ;
  LAYER metal2 ;
  RECT 615.440 763.280 618.980 764.400 ;
  LAYER metal1 ;
  RECT 615.440 763.280 618.980 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 572.040 763.280 575.580 764.400 ;
  LAYER metal3 ;
  RECT 572.040 763.280 575.580 764.400 ;
  LAYER metal2 ;
  RECT 572.040 763.280 575.580 764.400 ;
  LAYER metal1 ;
  RECT 572.040 763.280 575.580 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 563.360 763.280 566.900 764.400 ;
  LAYER metal3 ;
  RECT 563.360 763.280 566.900 764.400 ;
  LAYER metal2 ;
  RECT 563.360 763.280 566.900 764.400 ;
  LAYER metal1 ;
  RECT 563.360 763.280 566.900 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 554.680 763.280 558.220 764.400 ;
  LAYER metal3 ;
  RECT 554.680 763.280 558.220 764.400 ;
  LAYER metal2 ;
  RECT 554.680 763.280 558.220 764.400 ;
  LAYER metal1 ;
  RECT 554.680 763.280 558.220 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 546.000 763.280 549.540 764.400 ;
  LAYER metal3 ;
  RECT 546.000 763.280 549.540 764.400 ;
  LAYER metal2 ;
  RECT 546.000 763.280 549.540 764.400 ;
  LAYER metal1 ;
  RECT 546.000 763.280 549.540 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 537.320 763.280 540.860 764.400 ;
  LAYER metal3 ;
  RECT 537.320 763.280 540.860 764.400 ;
  LAYER metal2 ;
  RECT 537.320 763.280 540.860 764.400 ;
  LAYER metal1 ;
  RECT 537.320 763.280 540.860 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 528.640 763.280 532.180 764.400 ;
  LAYER metal3 ;
  RECT 528.640 763.280 532.180 764.400 ;
  LAYER metal2 ;
  RECT 528.640 763.280 532.180 764.400 ;
  LAYER metal1 ;
  RECT 528.640 763.280 532.180 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 485.240 763.280 488.780 764.400 ;
  LAYER metal3 ;
  RECT 485.240 763.280 488.780 764.400 ;
  LAYER metal2 ;
  RECT 485.240 763.280 488.780 764.400 ;
  LAYER metal1 ;
  RECT 485.240 763.280 488.780 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 476.560 763.280 480.100 764.400 ;
  LAYER metal3 ;
  RECT 476.560 763.280 480.100 764.400 ;
  LAYER metal2 ;
  RECT 476.560 763.280 480.100 764.400 ;
  LAYER metal1 ;
  RECT 476.560 763.280 480.100 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 467.880 763.280 471.420 764.400 ;
  LAYER metal3 ;
  RECT 467.880 763.280 471.420 764.400 ;
  LAYER metal2 ;
  RECT 467.880 763.280 471.420 764.400 ;
  LAYER metal1 ;
  RECT 467.880 763.280 471.420 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 459.200 763.280 462.740 764.400 ;
  LAYER metal3 ;
  RECT 459.200 763.280 462.740 764.400 ;
  LAYER metal2 ;
  RECT 459.200 763.280 462.740 764.400 ;
  LAYER metal1 ;
  RECT 459.200 763.280 462.740 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 450.520 763.280 454.060 764.400 ;
  LAYER metal3 ;
  RECT 450.520 763.280 454.060 764.400 ;
  LAYER metal2 ;
  RECT 450.520 763.280 454.060 764.400 ;
  LAYER metal1 ;
  RECT 450.520 763.280 454.060 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 441.840 763.280 445.380 764.400 ;
  LAYER metal3 ;
  RECT 441.840 763.280 445.380 764.400 ;
  LAYER metal2 ;
  RECT 441.840 763.280 445.380 764.400 ;
  LAYER metal1 ;
  RECT 441.840 763.280 445.380 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 398.440 763.280 401.980 764.400 ;
  LAYER metal3 ;
  RECT 398.440 763.280 401.980 764.400 ;
  LAYER metal2 ;
  RECT 398.440 763.280 401.980 764.400 ;
  LAYER metal1 ;
  RECT 398.440 763.280 401.980 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 389.760 763.280 393.300 764.400 ;
  LAYER metal3 ;
  RECT 389.760 763.280 393.300 764.400 ;
  LAYER metal2 ;
  RECT 389.760 763.280 393.300 764.400 ;
  LAYER metal1 ;
  RECT 389.760 763.280 393.300 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 381.080 763.280 384.620 764.400 ;
  LAYER metal3 ;
  RECT 381.080 763.280 384.620 764.400 ;
  LAYER metal2 ;
  RECT 381.080 763.280 384.620 764.400 ;
  LAYER metal1 ;
  RECT 381.080 763.280 384.620 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 372.400 763.280 375.940 764.400 ;
  LAYER metal3 ;
  RECT 372.400 763.280 375.940 764.400 ;
  LAYER metal2 ;
  RECT 372.400 763.280 375.940 764.400 ;
  LAYER metal1 ;
  RECT 372.400 763.280 375.940 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 363.720 763.280 367.260 764.400 ;
  LAYER metal3 ;
  RECT 363.720 763.280 367.260 764.400 ;
  LAYER metal2 ;
  RECT 363.720 763.280 367.260 764.400 ;
  LAYER metal1 ;
  RECT 363.720 763.280 367.260 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 355.040 763.280 358.580 764.400 ;
  LAYER metal3 ;
  RECT 355.040 763.280 358.580 764.400 ;
  LAYER metal2 ;
  RECT 355.040 763.280 358.580 764.400 ;
  LAYER metal1 ;
  RECT 355.040 763.280 358.580 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 311.640 763.280 315.180 764.400 ;
  LAYER metal3 ;
  RECT 311.640 763.280 315.180 764.400 ;
  LAYER metal2 ;
  RECT 311.640 763.280 315.180 764.400 ;
  LAYER metal1 ;
  RECT 311.640 763.280 315.180 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 302.960 763.280 306.500 764.400 ;
  LAYER metal3 ;
  RECT 302.960 763.280 306.500 764.400 ;
  LAYER metal2 ;
  RECT 302.960 763.280 306.500 764.400 ;
  LAYER metal1 ;
  RECT 302.960 763.280 306.500 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 294.280 763.280 297.820 764.400 ;
  LAYER metal3 ;
  RECT 294.280 763.280 297.820 764.400 ;
  LAYER metal2 ;
  RECT 294.280 763.280 297.820 764.400 ;
  LAYER metal1 ;
  RECT 294.280 763.280 297.820 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 285.600 763.280 289.140 764.400 ;
  LAYER metal3 ;
  RECT 285.600 763.280 289.140 764.400 ;
  LAYER metal2 ;
  RECT 285.600 763.280 289.140 764.400 ;
  LAYER metal1 ;
  RECT 285.600 763.280 289.140 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 276.920 763.280 280.460 764.400 ;
  LAYER metal3 ;
  RECT 276.920 763.280 280.460 764.400 ;
  LAYER metal2 ;
  RECT 276.920 763.280 280.460 764.400 ;
  LAYER metal1 ;
  RECT 276.920 763.280 280.460 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 268.240 763.280 271.780 764.400 ;
  LAYER metal3 ;
  RECT 268.240 763.280 271.780 764.400 ;
  LAYER metal2 ;
  RECT 268.240 763.280 271.780 764.400 ;
  LAYER metal1 ;
  RECT 268.240 763.280 271.780 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 224.840 763.280 228.380 764.400 ;
  LAYER metal3 ;
  RECT 224.840 763.280 228.380 764.400 ;
  LAYER metal2 ;
  RECT 224.840 763.280 228.380 764.400 ;
  LAYER metal1 ;
  RECT 224.840 763.280 228.380 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 216.160 763.280 219.700 764.400 ;
  LAYER metal3 ;
  RECT 216.160 763.280 219.700 764.400 ;
  LAYER metal2 ;
  RECT 216.160 763.280 219.700 764.400 ;
  LAYER metal1 ;
  RECT 216.160 763.280 219.700 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 207.480 763.280 211.020 764.400 ;
  LAYER metal3 ;
  RECT 207.480 763.280 211.020 764.400 ;
  LAYER metal2 ;
  RECT 207.480 763.280 211.020 764.400 ;
  LAYER metal1 ;
  RECT 207.480 763.280 211.020 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 198.800 763.280 202.340 764.400 ;
  LAYER metal3 ;
  RECT 198.800 763.280 202.340 764.400 ;
  LAYER metal2 ;
  RECT 198.800 763.280 202.340 764.400 ;
  LAYER metal1 ;
  RECT 198.800 763.280 202.340 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.120 763.280 193.660 764.400 ;
  LAYER metal3 ;
  RECT 190.120 763.280 193.660 764.400 ;
  LAYER metal2 ;
  RECT 190.120 763.280 193.660 764.400 ;
  LAYER metal1 ;
  RECT 190.120 763.280 193.660 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 181.440 763.280 184.980 764.400 ;
  LAYER metal3 ;
  RECT 181.440 763.280 184.980 764.400 ;
  LAYER metal2 ;
  RECT 181.440 763.280 184.980 764.400 ;
  LAYER metal1 ;
  RECT 181.440 763.280 184.980 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 138.040 763.280 141.580 764.400 ;
  LAYER metal3 ;
  RECT 138.040 763.280 141.580 764.400 ;
  LAYER metal2 ;
  RECT 138.040 763.280 141.580 764.400 ;
  LAYER metal1 ;
  RECT 138.040 763.280 141.580 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 129.360 763.280 132.900 764.400 ;
  LAYER metal3 ;
  RECT 129.360 763.280 132.900 764.400 ;
  LAYER metal2 ;
  RECT 129.360 763.280 132.900 764.400 ;
  LAYER metal1 ;
  RECT 129.360 763.280 132.900 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 120.680 763.280 124.220 764.400 ;
  LAYER metal3 ;
  RECT 120.680 763.280 124.220 764.400 ;
  LAYER metal2 ;
  RECT 120.680 763.280 124.220 764.400 ;
  LAYER metal1 ;
  RECT 120.680 763.280 124.220 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 112.000 763.280 115.540 764.400 ;
  LAYER metal3 ;
  RECT 112.000 763.280 115.540 764.400 ;
  LAYER metal2 ;
  RECT 112.000 763.280 115.540 764.400 ;
  LAYER metal1 ;
  RECT 112.000 763.280 115.540 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 103.320 763.280 106.860 764.400 ;
  LAYER metal3 ;
  RECT 103.320 763.280 106.860 764.400 ;
  LAYER metal2 ;
  RECT 103.320 763.280 106.860 764.400 ;
  LAYER metal1 ;
  RECT 103.320 763.280 106.860 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 94.640 763.280 98.180 764.400 ;
  LAYER metal3 ;
  RECT 94.640 763.280 98.180 764.400 ;
  LAYER metal2 ;
  RECT 94.640 763.280 98.180 764.400 ;
  LAYER metal1 ;
  RECT 94.640 763.280 98.180 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 51.240 763.280 54.780 764.400 ;
  LAYER metal3 ;
  RECT 51.240 763.280 54.780 764.400 ;
  LAYER metal2 ;
  RECT 51.240 763.280 54.780 764.400 ;
  LAYER metal1 ;
  RECT 51.240 763.280 54.780 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 42.560 763.280 46.100 764.400 ;
  LAYER metal3 ;
  RECT 42.560 763.280 46.100 764.400 ;
  LAYER metal2 ;
  RECT 42.560 763.280 46.100 764.400 ;
  LAYER metal1 ;
  RECT 42.560 763.280 46.100 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 33.880 763.280 37.420 764.400 ;
  LAYER metal3 ;
  RECT 33.880 763.280 37.420 764.400 ;
  LAYER metal2 ;
  RECT 33.880 763.280 37.420 764.400 ;
  LAYER metal1 ;
  RECT 33.880 763.280 37.420 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.200 763.280 28.740 764.400 ;
  LAYER metal3 ;
  RECT 25.200 763.280 28.740 764.400 ;
  LAYER metal2 ;
  RECT 25.200 763.280 28.740 764.400 ;
  LAYER metal1 ;
  RECT 25.200 763.280 28.740 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 16.520 763.280 20.060 764.400 ;
  LAYER metal3 ;
  RECT 16.520 763.280 20.060 764.400 ;
  LAYER metal2 ;
  RECT 16.520 763.280 20.060 764.400 ;
  LAYER metal1 ;
  RECT 16.520 763.280 20.060 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.840 763.280 11.380 764.400 ;
  LAYER metal3 ;
  RECT 7.840 763.280 11.380 764.400 ;
  LAYER metal2 ;
  RECT 7.840 763.280 11.380 764.400 ;
  LAYER metal1 ;
  RECT 7.840 763.280 11.380 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1004.180 0.000 1007.720 1.120 ;
  LAYER metal3 ;
  RECT 1004.180 0.000 1007.720 1.120 ;
  LAYER metal2 ;
  RECT 1004.180 0.000 1007.720 1.120 ;
  LAYER metal1 ;
  RECT 1004.180 0.000 1007.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 960.780 0.000 964.320 1.120 ;
  LAYER metal3 ;
  RECT 960.780 0.000 964.320 1.120 ;
  LAYER metal2 ;
  RECT 960.780 0.000 964.320 1.120 ;
  LAYER metal1 ;
  RECT 960.780 0.000 964.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 952.100 0.000 955.640 1.120 ;
  LAYER metal3 ;
  RECT 952.100 0.000 955.640 1.120 ;
  LAYER metal2 ;
  RECT 952.100 0.000 955.640 1.120 ;
  LAYER metal1 ;
  RECT 952.100 0.000 955.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 943.420 0.000 946.960 1.120 ;
  LAYER metal3 ;
  RECT 943.420 0.000 946.960 1.120 ;
  LAYER metal2 ;
  RECT 943.420 0.000 946.960 1.120 ;
  LAYER metal1 ;
  RECT 943.420 0.000 946.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 934.740 0.000 938.280 1.120 ;
  LAYER metal3 ;
  RECT 934.740 0.000 938.280 1.120 ;
  LAYER metal2 ;
  RECT 934.740 0.000 938.280 1.120 ;
  LAYER metal1 ;
  RECT 934.740 0.000 938.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 926.060 0.000 929.600 1.120 ;
  LAYER metal3 ;
  RECT 926.060 0.000 929.600 1.120 ;
  LAYER metal2 ;
  RECT 926.060 0.000 929.600 1.120 ;
  LAYER metal1 ;
  RECT 926.060 0.000 929.600 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 917.380 0.000 920.920 1.120 ;
  LAYER metal3 ;
  RECT 917.380 0.000 920.920 1.120 ;
  LAYER metal2 ;
  RECT 917.380 0.000 920.920 1.120 ;
  LAYER metal1 ;
  RECT 917.380 0.000 920.920 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 873.980 0.000 877.520 1.120 ;
  LAYER metal3 ;
  RECT 873.980 0.000 877.520 1.120 ;
  LAYER metal2 ;
  RECT 873.980 0.000 877.520 1.120 ;
  LAYER metal1 ;
  RECT 873.980 0.000 877.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 865.300 0.000 868.840 1.120 ;
  LAYER metal3 ;
  RECT 865.300 0.000 868.840 1.120 ;
  LAYER metal2 ;
  RECT 865.300 0.000 868.840 1.120 ;
  LAYER metal1 ;
  RECT 865.300 0.000 868.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 856.620 0.000 860.160 1.120 ;
  LAYER metal3 ;
  RECT 856.620 0.000 860.160 1.120 ;
  LAYER metal2 ;
  RECT 856.620 0.000 860.160 1.120 ;
  LAYER metal1 ;
  RECT 856.620 0.000 860.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal3 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal2 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal1 ;
  RECT 847.940 0.000 851.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal3 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal2 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal1 ;
  RECT 839.260 0.000 842.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 830.580 0.000 834.120 1.120 ;
  LAYER metal3 ;
  RECT 830.580 0.000 834.120 1.120 ;
  LAYER metal2 ;
  RECT 830.580 0.000 834.120 1.120 ;
  LAYER metal1 ;
  RECT 830.580 0.000 834.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 769.820 0.000 773.360 1.120 ;
  LAYER metal3 ;
  RECT 769.820 0.000 773.360 1.120 ;
  LAYER metal2 ;
  RECT 769.820 0.000 773.360 1.120 ;
  LAYER metal1 ;
  RECT 769.820 0.000 773.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 761.140 0.000 764.680 1.120 ;
  LAYER metal3 ;
  RECT 761.140 0.000 764.680 1.120 ;
  LAYER metal2 ;
  RECT 761.140 0.000 764.680 1.120 ;
  LAYER metal1 ;
  RECT 761.140 0.000 764.680 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 752.460 0.000 756.000 1.120 ;
  LAYER metal3 ;
  RECT 752.460 0.000 756.000 1.120 ;
  LAYER metal2 ;
  RECT 752.460 0.000 756.000 1.120 ;
  LAYER metal1 ;
  RECT 752.460 0.000 756.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 743.780 0.000 747.320 1.120 ;
  LAYER metal3 ;
  RECT 743.780 0.000 747.320 1.120 ;
  LAYER metal2 ;
  RECT 743.780 0.000 747.320 1.120 ;
  LAYER metal1 ;
  RECT 743.780 0.000 747.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 735.100 0.000 738.640 1.120 ;
  LAYER metal3 ;
  RECT 735.100 0.000 738.640 1.120 ;
  LAYER metal2 ;
  RECT 735.100 0.000 738.640 1.120 ;
  LAYER metal1 ;
  RECT 735.100 0.000 738.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 726.420 0.000 729.960 1.120 ;
  LAYER metal3 ;
  RECT 726.420 0.000 729.960 1.120 ;
  LAYER metal2 ;
  RECT 726.420 0.000 729.960 1.120 ;
  LAYER metal1 ;
  RECT 726.420 0.000 729.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 683.020 0.000 686.560 1.120 ;
  LAYER metal3 ;
  RECT 683.020 0.000 686.560 1.120 ;
  LAYER metal2 ;
  RECT 683.020 0.000 686.560 1.120 ;
  LAYER metal1 ;
  RECT 683.020 0.000 686.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 674.340 0.000 677.880 1.120 ;
  LAYER metal3 ;
  RECT 674.340 0.000 677.880 1.120 ;
  LAYER metal2 ;
  RECT 674.340 0.000 677.880 1.120 ;
  LAYER metal1 ;
  RECT 674.340 0.000 677.880 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 665.660 0.000 669.200 1.120 ;
  LAYER metal3 ;
  RECT 665.660 0.000 669.200 1.120 ;
  LAYER metal2 ;
  RECT 665.660 0.000 669.200 1.120 ;
  LAYER metal1 ;
  RECT 665.660 0.000 669.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 656.980 0.000 660.520 1.120 ;
  LAYER metal3 ;
  RECT 656.980 0.000 660.520 1.120 ;
  LAYER metal2 ;
  RECT 656.980 0.000 660.520 1.120 ;
  LAYER metal1 ;
  RECT 656.980 0.000 660.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 648.300 0.000 651.840 1.120 ;
  LAYER metal3 ;
  RECT 648.300 0.000 651.840 1.120 ;
  LAYER metal2 ;
  RECT 648.300 0.000 651.840 1.120 ;
  LAYER metal1 ;
  RECT 648.300 0.000 651.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 639.620 0.000 643.160 1.120 ;
  LAYER metal3 ;
  RECT 639.620 0.000 643.160 1.120 ;
  LAYER metal2 ;
  RECT 639.620 0.000 643.160 1.120 ;
  LAYER metal1 ;
  RECT 639.620 0.000 643.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER metal3 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER metal2 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER metal1 ;
  RECT 596.220 0.000 599.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 587.540 0.000 591.080 1.120 ;
  LAYER metal3 ;
  RECT 587.540 0.000 591.080 1.120 ;
  LAYER metal2 ;
  RECT 587.540 0.000 591.080 1.120 ;
  LAYER metal1 ;
  RECT 587.540 0.000 591.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER metal3 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER metal2 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER metal1 ;
  RECT 578.860 0.000 582.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal3 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal2 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal1 ;
  RECT 557.160 0.000 560.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 521.200 0.000 524.740 1.120 ;
  LAYER metal3 ;
  RECT 521.200 0.000 524.740 1.120 ;
  LAYER metal2 ;
  RECT 521.200 0.000 524.740 1.120 ;
  LAYER metal1 ;
  RECT 521.200 0.000 524.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 493.300 0.000 496.840 1.120 ;
  LAYER metal3 ;
  RECT 493.300 0.000 496.840 1.120 ;
  LAYER metal2 ;
  RECT 493.300 0.000 496.840 1.120 ;
  LAYER metal1 ;
  RECT 493.300 0.000 496.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 435.020 0.000 438.560 1.120 ;
  LAYER metal3 ;
  RECT 435.020 0.000 438.560 1.120 ;
  LAYER metal2 ;
  RECT 435.020 0.000 438.560 1.120 ;
  LAYER metal1 ;
  RECT 435.020 0.000 438.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 426.340 0.000 429.880 1.120 ;
  LAYER metal3 ;
  RECT 426.340 0.000 429.880 1.120 ;
  LAYER metal2 ;
  RECT 426.340 0.000 429.880 1.120 ;
  LAYER metal1 ;
  RECT 426.340 0.000 429.880 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 417.660 0.000 421.200 1.120 ;
  LAYER metal3 ;
  RECT 417.660 0.000 421.200 1.120 ;
  LAYER metal2 ;
  RECT 417.660 0.000 421.200 1.120 ;
  LAYER metal1 ;
  RECT 417.660 0.000 421.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal3 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal2 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal1 ;
  RECT 408.980 0.000 412.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 400.300 0.000 403.840 1.120 ;
  LAYER metal3 ;
  RECT 400.300 0.000 403.840 1.120 ;
  LAYER metal2 ;
  RECT 400.300 0.000 403.840 1.120 ;
  LAYER metal1 ;
  RECT 400.300 0.000 403.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 391.620 0.000 395.160 1.120 ;
  LAYER metal3 ;
  RECT 391.620 0.000 395.160 1.120 ;
  LAYER metal2 ;
  RECT 391.620 0.000 395.160 1.120 ;
  LAYER metal1 ;
  RECT 391.620 0.000 395.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 348.220 0.000 351.760 1.120 ;
  LAYER metal3 ;
  RECT 348.220 0.000 351.760 1.120 ;
  LAYER metal2 ;
  RECT 348.220 0.000 351.760 1.120 ;
  LAYER metal1 ;
  RECT 348.220 0.000 351.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal3 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal2 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal1 ;
  RECT 339.540 0.000 343.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER metal3 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER metal2 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER metal1 ;
  RECT 330.860 0.000 334.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 322.180 0.000 325.720 1.120 ;
  LAYER metal3 ;
  RECT 322.180 0.000 325.720 1.120 ;
  LAYER metal2 ;
  RECT 322.180 0.000 325.720 1.120 ;
  LAYER metal1 ;
  RECT 322.180 0.000 325.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 313.500 0.000 317.040 1.120 ;
  LAYER metal3 ;
  RECT 313.500 0.000 317.040 1.120 ;
  LAYER metal2 ;
  RECT 313.500 0.000 317.040 1.120 ;
  LAYER metal1 ;
  RECT 313.500 0.000 317.040 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 304.820 0.000 308.360 1.120 ;
  LAYER metal3 ;
  RECT 304.820 0.000 308.360 1.120 ;
  LAYER metal2 ;
  RECT 304.820 0.000 308.360 1.120 ;
  LAYER metal1 ;
  RECT 304.820 0.000 308.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal3 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal2 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal1 ;
  RECT 261.420 0.000 264.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal3 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal2 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal1 ;
  RECT 239.720 0.000 243.260 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 226.700 0.000 230.240 1.120 ;
  LAYER metal3 ;
  RECT 226.700 0.000 230.240 1.120 ;
  LAYER metal2 ;
  RECT 226.700 0.000 230.240 1.120 ;
  LAYER metal1 ;
  RECT 226.700 0.000 230.240 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 218.020 0.000 221.560 1.120 ;
  LAYER metal3 ;
  RECT 218.020 0.000 221.560 1.120 ;
  LAYER metal2 ;
  RECT 218.020 0.000 221.560 1.120 ;
  LAYER metal1 ;
  RECT 218.020 0.000 221.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 209.340 0.000 212.880 1.120 ;
  LAYER metal3 ;
  RECT 209.340 0.000 212.880 1.120 ;
  LAYER metal2 ;
  RECT 209.340 0.000 212.880 1.120 ;
  LAYER metal1 ;
  RECT 209.340 0.000 212.880 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 200.660 0.000 204.200 1.120 ;
  LAYER metal3 ;
  RECT 200.660 0.000 204.200 1.120 ;
  LAYER metal2 ;
  RECT 200.660 0.000 204.200 1.120 ;
  LAYER metal1 ;
  RECT 200.660 0.000 204.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 157.260 0.000 160.800 1.120 ;
  LAYER metal3 ;
  RECT 157.260 0.000 160.800 1.120 ;
  LAYER metal2 ;
  RECT 157.260 0.000 160.800 1.120 ;
  LAYER metal1 ;
  RECT 157.260 0.000 160.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER metal3 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER metal2 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER metal1 ;
  RECT 148.580 0.000 152.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 131.220 0.000 134.760 1.120 ;
  LAYER metal3 ;
  RECT 131.220 0.000 134.760 1.120 ;
  LAYER metal2 ;
  RECT 131.220 0.000 134.760 1.120 ;
  LAYER metal1 ;
  RECT 131.220 0.000 134.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 122.540 0.000 126.080 1.120 ;
  LAYER metal3 ;
  RECT 122.540 0.000 126.080 1.120 ;
  LAYER metal2 ;
  RECT 122.540 0.000 126.080 1.120 ;
  LAYER metal1 ;
  RECT 122.540 0.000 126.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER metal3 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER metal2 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER metal1 ;
  RECT 61.780 0.000 65.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER metal3 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER metal2 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER metal1 ;
  RECT 53.100 0.000 56.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER metal3 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER metal2 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER metal1 ;
  RECT 44.420 0.000 47.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 1014.440 749.060 1015.560 752.300 ;
  LAYER metal3 ;
  RECT 1014.440 749.060 1015.560 752.300 ;
  LAYER metal2 ;
  RECT 1014.440 749.060 1015.560 752.300 ;
  LAYER metal1 ;
  RECT 1014.440 749.060 1015.560 752.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 741.220 1015.560 744.460 ;
  LAYER metal3 ;
  RECT 1014.440 741.220 1015.560 744.460 ;
  LAYER metal2 ;
  RECT 1014.440 741.220 1015.560 744.460 ;
  LAYER metal1 ;
  RECT 1014.440 741.220 1015.560 744.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 733.380 1015.560 736.620 ;
  LAYER metal3 ;
  RECT 1014.440 733.380 1015.560 736.620 ;
  LAYER metal2 ;
  RECT 1014.440 733.380 1015.560 736.620 ;
  LAYER metal1 ;
  RECT 1014.440 733.380 1015.560 736.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 725.540 1015.560 728.780 ;
  LAYER metal3 ;
  RECT 1014.440 725.540 1015.560 728.780 ;
  LAYER metal2 ;
  RECT 1014.440 725.540 1015.560 728.780 ;
  LAYER metal1 ;
  RECT 1014.440 725.540 1015.560 728.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 717.700 1015.560 720.940 ;
  LAYER metal3 ;
  RECT 1014.440 717.700 1015.560 720.940 ;
  LAYER metal2 ;
  RECT 1014.440 717.700 1015.560 720.940 ;
  LAYER metal1 ;
  RECT 1014.440 717.700 1015.560 720.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 678.500 1015.560 681.740 ;
  LAYER metal3 ;
  RECT 1014.440 678.500 1015.560 681.740 ;
  LAYER metal2 ;
  RECT 1014.440 678.500 1015.560 681.740 ;
  LAYER metal1 ;
  RECT 1014.440 678.500 1015.560 681.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 670.660 1015.560 673.900 ;
  LAYER metal3 ;
  RECT 1014.440 670.660 1015.560 673.900 ;
  LAYER metal2 ;
  RECT 1014.440 670.660 1015.560 673.900 ;
  LAYER metal1 ;
  RECT 1014.440 670.660 1015.560 673.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 662.820 1015.560 666.060 ;
  LAYER metal3 ;
  RECT 1014.440 662.820 1015.560 666.060 ;
  LAYER metal2 ;
  RECT 1014.440 662.820 1015.560 666.060 ;
  LAYER metal1 ;
  RECT 1014.440 662.820 1015.560 666.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 654.980 1015.560 658.220 ;
  LAYER metal3 ;
  RECT 1014.440 654.980 1015.560 658.220 ;
  LAYER metal2 ;
  RECT 1014.440 654.980 1015.560 658.220 ;
  LAYER metal1 ;
  RECT 1014.440 654.980 1015.560 658.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 647.140 1015.560 650.380 ;
  LAYER metal3 ;
  RECT 1014.440 647.140 1015.560 650.380 ;
  LAYER metal2 ;
  RECT 1014.440 647.140 1015.560 650.380 ;
  LAYER metal1 ;
  RECT 1014.440 647.140 1015.560 650.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 639.300 1015.560 642.540 ;
  LAYER metal3 ;
  RECT 1014.440 639.300 1015.560 642.540 ;
  LAYER metal2 ;
  RECT 1014.440 639.300 1015.560 642.540 ;
  LAYER metal1 ;
  RECT 1014.440 639.300 1015.560 642.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 600.100 1015.560 603.340 ;
  LAYER metal3 ;
  RECT 1014.440 600.100 1015.560 603.340 ;
  LAYER metal2 ;
  RECT 1014.440 600.100 1015.560 603.340 ;
  LAYER metal1 ;
  RECT 1014.440 600.100 1015.560 603.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 592.260 1015.560 595.500 ;
  LAYER metal3 ;
  RECT 1014.440 592.260 1015.560 595.500 ;
  LAYER metal2 ;
  RECT 1014.440 592.260 1015.560 595.500 ;
  LAYER metal1 ;
  RECT 1014.440 592.260 1015.560 595.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 584.420 1015.560 587.660 ;
  LAYER metal3 ;
  RECT 1014.440 584.420 1015.560 587.660 ;
  LAYER metal2 ;
  RECT 1014.440 584.420 1015.560 587.660 ;
  LAYER metal1 ;
  RECT 1014.440 584.420 1015.560 587.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 576.580 1015.560 579.820 ;
  LAYER metal3 ;
  RECT 1014.440 576.580 1015.560 579.820 ;
  LAYER metal2 ;
  RECT 1014.440 576.580 1015.560 579.820 ;
  LAYER metal1 ;
  RECT 1014.440 576.580 1015.560 579.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 568.740 1015.560 571.980 ;
  LAYER metal3 ;
  RECT 1014.440 568.740 1015.560 571.980 ;
  LAYER metal2 ;
  RECT 1014.440 568.740 1015.560 571.980 ;
  LAYER metal1 ;
  RECT 1014.440 568.740 1015.560 571.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 560.900 1015.560 564.140 ;
  LAYER metal3 ;
  RECT 1014.440 560.900 1015.560 564.140 ;
  LAYER metal2 ;
  RECT 1014.440 560.900 1015.560 564.140 ;
  LAYER metal1 ;
  RECT 1014.440 560.900 1015.560 564.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 521.700 1015.560 524.940 ;
  LAYER metal3 ;
  RECT 1014.440 521.700 1015.560 524.940 ;
  LAYER metal2 ;
  RECT 1014.440 521.700 1015.560 524.940 ;
  LAYER metal1 ;
  RECT 1014.440 521.700 1015.560 524.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 513.860 1015.560 517.100 ;
  LAYER metal3 ;
  RECT 1014.440 513.860 1015.560 517.100 ;
  LAYER metal2 ;
  RECT 1014.440 513.860 1015.560 517.100 ;
  LAYER metal1 ;
  RECT 1014.440 513.860 1015.560 517.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 506.020 1015.560 509.260 ;
  LAYER metal3 ;
  RECT 1014.440 506.020 1015.560 509.260 ;
  LAYER metal2 ;
  RECT 1014.440 506.020 1015.560 509.260 ;
  LAYER metal1 ;
  RECT 1014.440 506.020 1015.560 509.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 498.180 1015.560 501.420 ;
  LAYER metal3 ;
  RECT 1014.440 498.180 1015.560 501.420 ;
  LAYER metal2 ;
  RECT 1014.440 498.180 1015.560 501.420 ;
  LAYER metal1 ;
  RECT 1014.440 498.180 1015.560 501.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 490.340 1015.560 493.580 ;
  LAYER metal3 ;
  RECT 1014.440 490.340 1015.560 493.580 ;
  LAYER metal2 ;
  RECT 1014.440 490.340 1015.560 493.580 ;
  LAYER metal1 ;
  RECT 1014.440 490.340 1015.560 493.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 482.500 1015.560 485.740 ;
  LAYER metal3 ;
  RECT 1014.440 482.500 1015.560 485.740 ;
  LAYER metal2 ;
  RECT 1014.440 482.500 1015.560 485.740 ;
  LAYER metal1 ;
  RECT 1014.440 482.500 1015.560 485.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 443.300 1015.560 446.540 ;
  LAYER metal3 ;
  RECT 1014.440 443.300 1015.560 446.540 ;
  LAYER metal2 ;
  RECT 1014.440 443.300 1015.560 446.540 ;
  LAYER metal1 ;
  RECT 1014.440 443.300 1015.560 446.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 435.460 1015.560 438.700 ;
  LAYER metal3 ;
  RECT 1014.440 435.460 1015.560 438.700 ;
  LAYER metal2 ;
  RECT 1014.440 435.460 1015.560 438.700 ;
  LAYER metal1 ;
  RECT 1014.440 435.460 1015.560 438.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 427.620 1015.560 430.860 ;
  LAYER metal3 ;
  RECT 1014.440 427.620 1015.560 430.860 ;
  LAYER metal2 ;
  RECT 1014.440 427.620 1015.560 430.860 ;
  LAYER metal1 ;
  RECT 1014.440 427.620 1015.560 430.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 419.780 1015.560 423.020 ;
  LAYER metal3 ;
  RECT 1014.440 419.780 1015.560 423.020 ;
  LAYER metal2 ;
  RECT 1014.440 419.780 1015.560 423.020 ;
  LAYER metal1 ;
  RECT 1014.440 419.780 1015.560 423.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 411.940 1015.560 415.180 ;
  LAYER metal3 ;
  RECT 1014.440 411.940 1015.560 415.180 ;
  LAYER metal2 ;
  RECT 1014.440 411.940 1015.560 415.180 ;
  LAYER metal1 ;
  RECT 1014.440 411.940 1015.560 415.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 404.100 1015.560 407.340 ;
  LAYER metal3 ;
  RECT 1014.440 404.100 1015.560 407.340 ;
  LAYER metal2 ;
  RECT 1014.440 404.100 1015.560 407.340 ;
  LAYER metal1 ;
  RECT 1014.440 404.100 1015.560 407.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 364.900 1015.560 368.140 ;
  LAYER metal3 ;
  RECT 1014.440 364.900 1015.560 368.140 ;
  LAYER metal2 ;
  RECT 1014.440 364.900 1015.560 368.140 ;
  LAYER metal1 ;
  RECT 1014.440 364.900 1015.560 368.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 357.060 1015.560 360.300 ;
  LAYER metal3 ;
  RECT 1014.440 357.060 1015.560 360.300 ;
  LAYER metal2 ;
  RECT 1014.440 357.060 1015.560 360.300 ;
  LAYER metal1 ;
  RECT 1014.440 357.060 1015.560 360.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 349.220 1015.560 352.460 ;
  LAYER metal3 ;
  RECT 1014.440 349.220 1015.560 352.460 ;
  LAYER metal2 ;
  RECT 1014.440 349.220 1015.560 352.460 ;
  LAYER metal1 ;
  RECT 1014.440 349.220 1015.560 352.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 341.380 1015.560 344.620 ;
  LAYER metal3 ;
  RECT 1014.440 341.380 1015.560 344.620 ;
  LAYER metal2 ;
  RECT 1014.440 341.380 1015.560 344.620 ;
  LAYER metal1 ;
  RECT 1014.440 341.380 1015.560 344.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 333.540 1015.560 336.780 ;
  LAYER metal3 ;
  RECT 1014.440 333.540 1015.560 336.780 ;
  LAYER metal2 ;
  RECT 1014.440 333.540 1015.560 336.780 ;
  LAYER metal1 ;
  RECT 1014.440 333.540 1015.560 336.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 325.700 1015.560 328.940 ;
  LAYER metal3 ;
  RECT 1014.440 325.700 1015.560 328.940 ;
  LAYER metal2 ;
  RECT 1014.440 325.700 1015.560 328.940 ;
  LAYER metal1 ;
  RECT 1014.440 325.700 1015.560 328.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 286.500 1015.560 289.740 ;
  LAYER metal3 ;
  RECT 1014.440 286.500 1015.560 289.740 ;
  LAYER metal2 ;
  RECT 1014.440 286.500 1015.560 289.740 ;
  LAYER metal1 ;
  RECT 1014.440 286.500 1015.560 289.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 278.660 1015.560 281.900 ;
  LAYER metal3 ;
  RECT 1014.440 278.660 1015.560 281.900 ;
  LAYER metal2 ;
  RECT 1014.440 278.660 1015.560 281.900 ;
  LAYER metal1 ;
  RECT 1014.440 278.660 1015.560 281.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 270.820 1015.560 274.060 ;
  LAYER metal3 ;
  RECT 1014.440 270.820 1015.560 274.060 ;
  LAYER metal2 ;
  RECT 1014.440 270.820 1015.560 274.060 ;
  LAYER metal1 ;
  RECT 1014.440 270.820 1015.560 274.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 262.980 1015.560 266.220 ;
  LAYER metal3 ;
  RECT 1014.440 262.980 1015.560 266.220 ;
  LAYER metal2 ;
  RECT 1014.440 262.980 1015.560 266.220 ;
  LAYER metal1 ;
  RECT 1014.440 262.980 1015.560 266.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 255.140 1015.560 258.380 ;
  LAYER metal3 ;
  RECT 1014.440 255.140 1015.560 258.380 ;
  LAYER metal2 ;
  RECT 1014.440 255.140 1015.560 258.380 ;
  LAYER metal1 ;
  RECT 1014.440 255.140 1015.560 258.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 247.300 1015.560 250.540 ;
  LAYER metal3 ;
  RECT 1014.440 247.300 1015.560 250.540 ;
  LAYER metal2 ;
  RECT 1014.440 247.300 1015.560 250.540 ;
  LAYER metal1 ;
  RECT 1014.440 247.300 1015.560 250.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 208.100 1015.560 211.340 ;
  LAYER metal3 ;
  RECT 1014.440 208.100 1015.560 211.340 ;
  LAYER metal2 ;
  RECT 1014.440 208.100 1015.560 211.340 ;
  LAYER metal1 ;
  RECT 1014.440 208.100 1015.560 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 200.260 1015.560 203.500 ;
  LAYER metal3 ;
  RECT 1014.440 200.260 1015.560 203.500 ;
  LAYER metal2 ;
  RECT 1014.440 200.260 1015.560 203.500 ;
  LAYER metal1 ;
  RECT 1014.440 200.260 1015.560 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 192.420 1015.560 195.660 ;
  LAYER metal3 ;
  RECT 1014.440 192.420 1015.560 195.660 ;
  LAYER metal2 ;
  RECT 1014.440 192.420 1015.560 195.660 ;
  LAYER metal1 ;
  RECT 1014.440 192.420 1015.560 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 184.580 1015.560 187.820 ;
  LAYER metal3 ;
  RECT 1014.440 184.580 1015.560 187.820 ;
  LAYER metal2 ;
  RECT 1014.440 184.580 1015.560 187.820 ;
  LAYER metal1 ;
  RECT 1014.440 184.580 1015.560 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 176.740 1015.560 179.980 ;
  LAYER metal3 ;
  RECT 1014.440 176.740 1015.560 179.980 ;
  LAYER metal2 ;
  RECT 1014.440 176.740 1015.560 179.980 ;
  LAYER metal1 ;
  RECT 1014.440 176.740 1015.560 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 168.900 1015.560 172.140 ;
  LAYER metal3 ;
  RECT 1014.440 168.900 1015.560 172.140 ;
  LAYER metal2 ;
  RECT 1014.440 168.900 1015.560 172.140 ;
  LAYER metal1 ;
  RECT 1014.440 168.900 1015.560 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 129.700 1015.560 132.940 ;
  LAYER metal3 ;
  RECT 1014.440 129.700 1015.560 132.940 ;
  LAYER metal2 ;
  RECT 1014.440 129.700 1015.560 132.940 ;
  LAYER metal1 ;
  RECT 1014.440 129.700 1015.560 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 121.860 1015.560 125.100 ;
  LAYER metal3 ;
  RECT 1014.440 121.860 1015.560 125.100 ;
  LAYER metal2 ;
  RECT 1014.440 121.860 1015.560 125.100 ;
  LAYER metal1 ;
  RECT 1014.440 121.860 1015.560 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 114.020 1015.560 117.260 ;
  LAYER metal3 ;
  RECT 1014.440 114.020 1015.560 117.260 ;
  LAYER metal2 ;
  RECT 1014.440 114.020 1015.560 117.260 ;
  LAYER metal1 ;
  RECT 1014.440 114.020 1015.560 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 106.180 1015.560 109.420 ;
  LAYER metal3 ;
  RECT 1014.440 106.180 1015.560 109.420 ;
  LAYER metal2 ;
  RECT 1014.440 106.180 1015.560 109.420 ;
  LAYER metal1 ;
  RECT 1014.440 106.180 1015.560 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 98.340 1015.560 101.580 ;
  LAYER metal3 ;
  RECT 1014.440 98.340 1015.560 101.580 ;
  LAYER metal2 ;
  RECT 1014.440 98.340 1015.560 101.580 ;
  LAYER metal1 ;
  RECT 1014.440 98.340 1015.560 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 90.500 1015.560 93.740 ;
  LAYER metal3 ;
  RECT 1014.440 90.500 1015.560 93.740 ;
  LAYER metal2 ;
  RECT 1014.440 90.500 1015.560 93.740 ;
  LAYER metal1 ;
  RECT 1014.440 90.500 1015.560 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 51.300 1015.560 54.540 ;
  LAYER metal3 ;
  RECT 1014.440 51.300 1015.560 54.540 ;
  LAYER metal2 ;
  RECT 1014.440 51.300 1015.560 54.540 ;
  LAYER metal1 ;
  RECT 1014.440 51.300 1015.560 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 43.460 1015.560 46.700 ;
  LAYER metal3 ;
  RECT 1014.440 43.460 1015.560 46.700 ;
  LAYER metal2 ;
  RECT 1014.440 43.460 1015.560 46.700 ;
  LAYER metal1 ;
  RECT 1014.440 43.460 1015.560 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 35.620 1015.560 38.860 ;
  LAYER metal3 ;
  RECT 1014.440 35.620 1015.560 38.860 ;
  LAYER metal2 ;
  RECT 1014.440 35.620 1015.560 38.860 ;
  LAYER metal1 ;
  RECT 1014.440 35.620 1015.560 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 27.780 1015.560 31.020 ;
  LAYER metal3 ;
  RECT 1014.440 27.780 1015.560 31.020 ;
  LAYER metal2 ;
  RECT 1014.440 27.780 1015.560 31.020 ;
  LAYER metal1 ;
  RECT 1014.440 27.780 1015.560 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 19.940 1015.560 23.180 ;
  LAYER metal3 ;
  RECT 1014.440 19.940 1015.560 23.180 ;
  LAYER metal2 ;
  RECT 1014.440 19.940 1015.560 23.180 ;
  LAYER metal1 ;
  RECT 1014.440 19.940 1015.560 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.440 12.100 1015.560 15.340 ;
  LAYER metal3 ;
  RECT 1014.440 12.100 1015.560 15.340 ;
  LAYER metal2 ;
  RECT 1014.440 12.100 1015.560 15.340 ;
  LAYER metal1 ;
  RECT 1014.440 12.100 1015.560 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 749.060 1.120 752.300 ;
  LAYER metal3 ;
  RECT 0.000 749.060 1.120 752.300 ;
  LAYER metal2 ;
  RECT 0.000 749.060 1.120 752.300 ;
  LAYER metal1 ;
  RECT 0.000 749.060 1.120 752.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 741.220 1.120 744.460 ;
  LAYER metal3 ;
  RECT 0.000 741.220 1.120 744.460 ;
  LAYER metal2 ;
  RECT 0.000 741.220 1.120 744.460 ;
  LAYER metal1 ;
  RECT 0.000 741.220 1.120 744.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 733.380 1.120 736.620 ;
  LAYER metal3 ;
  RECT 0.000 733.380 1.120 736.620 ;
  LAYER metal2 ;
  RECT 0.000 733.380 1.120 736.620 ;
  LAYER metal1 ;
  RECT 0.000 733.380 1.120 736.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 725.540 1.120 728.780 ;
  LAYER metal3 ;
  RECT 0.000 725.540 1.120 728.780 ;
  LAYER metal2 ;
  RECT 0.000 725.540 1.120 728.780 ;
  LAYER metal1 ;
  RECT 0.000 725.540 1.120 728.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 717.700 1.120 720.940 ;
  LAYER metal3 ;
  RECT 0.000 717.700 1.120 720.940 ;
  LAYER metal2 ;
  RECT 0.000 717.700 1.120 720.940 ;
  LAYER metal1 ;
  RECT 0.000 717.700 1.120 720.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 678.500 1.120 681.740 ;
  LAYER metal3 ;
  RECT 0.000 678.500 1.120 681.740 ;
  LAYER metal2 ;
  RECT 0.000 678.500 1.120 681.740 ;
  LAYER metal1 ;
  RECT 0.000 678.500 1.120 681.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 670.660 1.120 673.900 ;
  LAYER metal3 ;
  RECT 0.000 670.660 1.120 673.900 ;
  LAYER metal2 ;
  RECT 0.000 670.660 1.120 673.900 ;
  LAYER metal1 ;
  RECT 0.000 670.660 1.120 673.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 662.820 1.120 666.060 ;
  LAYER metal3 ;
  RECT 0.000 662.820 1.120 666.060 ;
  LAYER metal2 ;
  RECT 0.000 662.820 1.120 666.060 ;
  LAYER metal1 ;
  RECT 0.000 662.820 1.120 666.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 654.980 1.120 658.220 ;
  LAYER metal3 ;
  RECT 0.000 654.980 1.120 658.220 ;
  LAYER metal2 ;
  RECT 0.000 654.980 1.120 658.220 ;
  LAYER metal1 ;
  RECT 0.000 654.980 1.120 658.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 647.140 1.120 650.380 ;
  LAYER metal3 ;
  RECT 0.000 647.140 1.120 650.380 ;
  LAYER metal2 ;
  RECT 0.000 647.140 1.120 650.380 ;
  LAYER metal1 ;
  RECT 0.000 647.140 1.120 650.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 639.300 1.120 642.540 ;
  LAYER metal3 ;
  RECT 0.000 639.300 1.120 642.540 ;
  LAYER metal2 ;
  RECT 0.000 639.300 1.120 642.540 ;
  LAYER metal1 ;
  RECT 0.000 639.300 1.120 642.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 600.100 1.120 603.340 ;
  LAYER metal3 ;
  RECT 0.000 600.100 1.120 603.340 ;
  LAYER metal2 ;
  RECT 0.000 600.100 1.120 603.340 ;
  LAYER metal1 ;
  RECT 0.000 600.100 1.120 603.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 592.260 1.120 595.500 ;
  LAYER metal3 ;
  RECT 0.000 592.260 1.120 595.500 ;
  LAYER metal2 ;
  RECT 0.000 592.260 1.120 595.500 ;
  LAYER metal1 ;
  RECT 0.000 592.260 1.120 595.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 584.420 1.120 587.660 ;
  LAYER metal3 ;
  RECT 0.000 584.420 1.120 587.660 ;
  LAYER metal2 ;
  RECT 0.000 584.420 1.120 587.660 ;
  LAYER metal1 ;
  RECT 0.000 584.420 1.120 587.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 576.580 1.120 579.820 ;
  LAYER metal3 ;
  RECT 0.000 576.580 1.120 579.820 ;
  LAYER metal2 ;
  RECT 0.000 576.580 1.120 579.820 ;
  LAYER metal1 ;
  RECT 0.000 576.580 1.120 579.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 568.740 1.120 571.980 ;
  LAYER metal3 ;
  RECT 0.000 568.740 1.120 571.980 ;
  LAYER metal2 ;
  RECT 0.000 568.740 1.120 571.980 ;
  LAYER metal1 ;
  RECT 0.000 568.740 1.120 571.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 560.900 1.120 564.140 ;
  LAYER metal3 ;
  RECT 0.000 560.900 1.120 564.140 ;
  LAYER metal2 ;
  RECT 0.000 560.900 1.120 564.140 ;
  LAYER metal1 ;
  RECT 0.000 560.900 1.120 564.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER metal3 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER metal2 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER metal1 ;
  RECT 0.000 521.700 1.120 524.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER metal3 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER metal2 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER metal1 ;
  RECT 0.000 513.860 1.120 517.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER metal3 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER metal2 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER metal1 ;
  RECT 0.000 506.020 1.120 509.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER metal3 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER metal2 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER metal1 ;
  RECT 0.000 498.180 1.120 501.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER metal3 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER metal2 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER metal1 ;
  RECT 0.000 490.340 1.120 493.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER metal3 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER metal2 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER metal1 ;
  RECT 0.000 482.500 1.120 485.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER metal3 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER metal2 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER metal1 ;
  RECT 0.000 443.300 1.120 446.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER metal3 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER metal2 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER metal1 ;
  RECT 0.000 435.460 1.120 438.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER metal3 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER metal2 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER metal1 ;
  RECT 0.000 427.620 1.120 430.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER metal3 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER metal2 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER metal1 ;
  RECT 0.000 419.780 1.120 423.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER metal3 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER metal2 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER metal1 ;
  RECT 0.000 411.940 1.120 415.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER metal3 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER metal2 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER metal1 ;
  RECT 0.000 404.100 1.120 407.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER metal3 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER metal2 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER metal1 ;
  RECT 0.000 364.900 1.120 368.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER metal3 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER metal2 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER metal1 ;
  RECT 0.000 357.060 1.120 360.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER metal3 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER metal2 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER metal1 ;
  RECT 0.000 349.220 1.120 352.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER metal3 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER metal2 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER metal1 ;
  RECT 0.000 341.380 1.120 344.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER metal3 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER metal2 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER metal1 ;
  RECT 0.000 333.540 1.120 336.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER metal3 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER metal2 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER metal1 ;
  RECT 0.000 325.700 1.120 328.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER metal3 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER metal2 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER metal1 ;
  RECT 0.000 286.500 1.120 289.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal3 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal2 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal1 ;
  RECT 0.000 278.660 1.120 281.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal3 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal2 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal1 ;
  RECT 0.000 270.820 1.120 274.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal3 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal2 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal1 ;
  RECT 0.000 262.980 1.120 266.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal3 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal2 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal1 ;
  RECT 0.000 255.140 1.120 258.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal3 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal2 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal1 ;
  RECT 0.000 247.300 1.120 250.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal3 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal2 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal1 ;
  RECT 0.000 208.100 1.120 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1001.700 763.280 1005.240 764.400 ;
  LAYER metal3 ;
  RECT 1001.700 763.280 1005.240 764.400 ;
  LAYER metal2 ;
  RECT 1001.700 763.280 1005.240 764.400 ;
  LAYER metal1 ;
  RECT 1001.700 763.280 1005.240 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 993.020 763.280 996.560 764.400 ;
  LAYER metal3 ;
  RECT 993.020 763.280 996.560 764.400 ;
  LAYER metal2 ;
  RECT 993.020 763.280 996.560 764.400 ;
  LAYER metal1 ;
  RECT 993.020 763.280 996.560 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 984.340 763.280 987.880 764.400 ;
  LAYER metal3 ;
  RECT 984.340 763.280 987.880 764.400 ;
  LAYER metal2 ;
  RECT 984.340 763.280 987.880 764.400 ;
  LAYER metal1 ;
  RECT 984.340 763.280 987.880 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 975.660 763.280 979.200 764.400 ;
  LAYER metal3 ;
  RECT 975.660 763.280 979.200 764.400 ;
  LAYER metal2 ;
  RECT 975.660 763.280 979.200 764.400 ;
  LAYER metal1 ;
  RECT 975.660 763.280 979.200 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 966.980 763.280 970.520 764.400 ;
  LAYER metal3 ;
  RECT 966.980 763.280 970.520 764.400 ;
  LAYER metal2 ;
  RECT 966.980 763.280 970.520 764.400 ;
  LAYER metal1 ;
  RECT 966.980 763.280 970.520 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 923.580 763.280 927.120 764.400 ;
  LAYER metal3 ;
  RECT 923.580 763.280 927.120 764.400 ;
  LAYER metal2 ;
  RECT 923.580 763.280 927.120 764.400 ;
  LAYER metal1 ;
  RECT 923.580 763.280 927.120 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 914.900 763.280 918.440 764.400 ;
  LAYER metal3 ;
  RECT 914.900 763.280 918.440 764.400 ;
  LAYER metal2 ;
  RECT 914.900 763.280 918.440 764.400 ;
  LAYER metal1 ;
  RECT 914.900 763.280 918.440 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 906.220 763.280 909.760 764.400 ;
  LAYER metal3 ;
  RECT 906.220 763.280 909.760 764.400 ;
  LAYER metal2 ;
  RECT 906.220 763.280 909.760 764.400 ;
  LAYER metal1 ;
  RECT 906.220 763.280 909.760 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 897.540 763.280 901.080 764.400 ;
  LAYER metal3 ;
  RECT 897.540 763.280 901.080 764.400 ;
  LAYER metal2 ;
  RECT 897.540 763.280 901.080 764.400 ;
  LAYER metal1 ;
  RECT 897.540 763.280 901.080 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 888.860 763.280 892.400 764.400 ;
  LAYER metal3 ;
  RECT 888.860 763.280 892.400 764.400 ;
  LAYER metal2 ;
  RECT 888.860 763.280 892.400 764.400 ;
  LAYER metal1 ;
  RECT 888.860 763.280 892.400 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 880.180 763.280 883.720 764.400 ;
  LAYER metal3 ;
  RECT 880.180 763.280 883.720 764.400 ;
  LAYER metal2 ;
  RECT 880.180 763.280 883.720 764.400 ;
  LAYER metal1 ;
  RECT 880.180 763.280 883.720 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 836.780 763.280 840.320 764.400 ;
  LAYER metal3 ;
  RECT 836.780 763.280 840.320 764.400 ;
  LAYER metal2 ;
  RECT 836.780 763.280 840.320 764.400 ;
  LAYER metal1 ;
  RECT 836.780 763.280 840.320 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 828.100 763.280 831.640 764.400 ;
  LAYER metal3 ;
  RECT 828.100 763.280 831.640 764.400 ;
  LAYER metal2 ;
  RECT 828.100 763.280 831.640 764.400 ;
  LAYER metal1 ;
  RECT 828.100 763.280 831.640 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 819.420 763.280 822.960 764.400 ;
  LAYER metal3 ;
  RECT 819.420 763.280 822.960 764.400 ;
  LAYER metal2 ;
  RECT 819.420 763.280 822.960 764.400 ;
  LAYER metal1 ;
  RECT 819.420 763.280 822.960 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 810.740 763.280 814.280 764.400 ;
  LAYER metal3 ;
  RECT 810.740 763.280 814.280 764.400 ;
  LAYER metal2 ;
  RECT 810.740 763.280 814.280 764.400 ;
  LAYER metal1 ;
  RECT 810.740 763.280 814.280 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 802.060 763.280 805.600 764.400 ;
  LAYER metal3 ;
  RECT 802.060 763.280 805.600 764.400 ;
  LAYER metal2 ;
  RECT 802.060 763.280 805.600 764.400 ;
  LAYER metal1 ;
  RECT 802.060 763.280 805.600 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 793.380 763.280 796.920 764.400 ;
  LAYER metal3 ;
  RECT 793.380 763.280 796.920 764.400 ;
  LAYER metal2 ;
  RECT 793.380 763.280 796.920 764.400 ;
  LAYER metal1 ;
  RECT 793.380 763.280 796.920 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.980 763.280 753.520 764.400 ;
  LAYER metal3 ;
  RECT 749.980 763.280 753.520 764.400 ;
  LAYER metal2 ;
  RECT 749.980 763.280 753.520 764.400 ;
  LAYER metal1 ;
  RECT 749.980 763.280 753.520 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 741.300 763.280 744.840 764.400 ;
  LAYER metal3 ;
  RECT 741.300 763.280 744.840 764.400 ;
  LAYER metal2 ;
  RECT 741.300 763.280 744.840 764.400 ;
  LAYER metal1 ;
  RECT 741.300 763.280 744.840 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 732.620 763.280 736.160 764.400 ;
  LAYER metal3 ;
  RECT 732.620 763.280 736.160 764.400 ;
  LAYER metal2 ;
  RECT 732.620 763.280 736.160 764.400 ;
  LAYER metal1 ;
  RECT 732.620 763.280 736.160 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 723.940 763.280 727.480 764.400 ;
  LAYER metal3 ;
  RECT 723.940 763.280 727.480 764.400 ;
  LAYER metal2 ;
  RECT 723.940 763.280 727.480 764.400 ;
  LAYER metal1 ;
  RECT 723.940 763.280 727.480 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 715.260 763.280 718.800 764.400 ;
  LAYER metal3 ;
  RECT 715.260 763.280 718.800 764.400 ;
  LAYER metal2 ;
  RECT 715.260 763.280 718.800 764.400 ;
  LAYER metal1 ;
  RECT 715.260 763.280 718.800 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 706.580 763.280 710.120 764.400 ;
  LAYER metal3 ;
  RECT 706.580 763.280 710.120 764.400 ;
  LAYER metal2 ;
  RECT 706.580 763.280 710.120 764.400 ;
  LAYER metal1 ;
  RECT 706.580 763.280 710.120 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 663.180 763.280 666.720 764.400 ;
  LAYER metal3 ;
  RECT 663.180 763.280 666.720 764.400 ;
  LAYER metal2 ;
  RECT 663.180 763.280 666.720 764.400 ;
  LAYER metal1 ;
  RECT 663.180 763.280 666.720 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 654.500 763.280 658.040 764.400 ;
  LAYER metal3 ;
  RECT 654.500 763.280 658.040 764.400 ;
  LAYER metal2 ;
  RECT 654.500 763.280 658.040 764.400 ;
  LAYER metal1 ;
  RECT 654.500 763.280 658.040 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 645.820 763.280 649.360 764.400 ;
  LAYER metal3 ;
  RECT 645.820 763.280 649.360 764.400 ;
  LAYER metal2 ;
  RECT 645.820 763.280 649.360 764.400 ;
  LAYER metal1 ;
  RECT 645.820 763.280 649.360 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 637.140 763.280 640.680 764.400 ;
  LAYER metal3 ;
  RECT 637.140 763.280 640.680 764.400 ;
  LAYER metal2 ;
  RECT 637.140 763.280 640.680 764.400 ;
  LAYER metal1 ;
  RECT 637.140 763.280 640.680 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 628.460 763.280 632.000 764.400 ;
  LAYER metal3 ;
  RECT 628.460 763.280 632.000 764.400 ;
  LAYER metal2 ;
  RECT 628.460 763.280 632.000 764.400 ;
  LAYER metal1 ;
  RECT 628.460 763.280 632.000 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 619.780 763.280 623.320 764.400 ;
  LAYER metal3 ;
  RECT 619.780 763.280 623.320 764.400 ;
  LAYER metal2 ;
  RECT 619.780 763.280 623.320 764.400 ;
  LAYER metal1 ;
  RECT 619.780 763.280 623.320 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 576.380 763.280 579.920 764.400 ;
  LAYER metal3 ;
  RECT 576.380 763.280 579.920 764.400 ;
  LAYER metal2 ;
  RECT 576.380 763.280 579.920 764.400 ;
  LAYER metal1 ;
  RECT 576.380 763.280 579.920 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 567.700 763.280 571.240 764.400 ;
  LAYER metal3 ;
  RECT 567.700 763.280 571.240 764.400 ;
  LAYER metal2 ;
  RECT 567.700 763.280 571.240 764.400 ;
  LAYER metal1 ;
  RECT 567.700 763.280 571.240 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 559.020 763.280 562.560 764.400 ;
  LAYER metal3 ;
  RECT 559.020 763.280 562.560 764.400 ;
  LAYER metal2 ;
  RECT 559.020 763.280 562.560 764.400 ;
  LAYER metal1 ;
  RECT 559.020 763.280 562.560 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 550.340 763.280 553.880 764.400 ;
  LAYER metal3 ;
  RECT 550.340 763.280 553.880 764.400 ;
  LAYER metal2 ;
  RECT 550.340 763.280 553.880 764.400 ;
  LAYER metal1 ;
  RECT 550.340 763.280 553.880 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 541.660 763.280 545.200 764.400 ;
  LAYER metal3 ;
  RECT 541.660 763.280 545.200 764.400 ;
  LAYER metal2 ;
  RECT 541.660 763.280 545.200 764.400 ;
  LAYER metal1 ;
  RECT 541.660 763.280 545.200 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 532.980 763.280 536.520 764.400 ;
  LAYER metal3 ;
  RECT 532.980 763.280 536.520 764.400 ;
  LAYER metal2 ;
  RECT 532.980 763.280 536.520 764.400 ;
  LAYER metal1 ;
  RECT 532.980 763.280 536.520 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 489.580 763.280 493.120 764.400 ;
  LAYER metal3 ;
  RECT 489.580 763.280 493.120 764.400 ;
  LAYER metal2 ;
  RECT 489.580 763.280 493.120 764.400 ;
  LAYER metal1 ;
  RECT 489.580 763.280 493.120 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 480.900 763.280 484.440 764.400 ;
  LAYER metal3 ;
  RECT 480.900 763.280 484.440 764.400 ;
  LAYER metal2 ;
  RECT 480.900 763.280 484.440 764.400 ;
  LAYER metal1 ;
  RECT 480.900 763.280 484.440 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 472.220 763.280 475.760 764.400 ;
  LAYER metal3 ;
  RECT 472.220 763.280 475.760 764.400 ;
  LAYER metal2 ;
  RECT 472.220 763.280 475.760 764.400 ;
  LAYER metal1 ;
  RECT 472.220 763.280 475.760 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 463.540 763.280 467.080 764.400 ;
  LAYER metal3 ;
  RECT 463.540 763.280 467.080 764.400 ;
  LAYER metal2 ;
  RECT 463.540 763.280 467.080 764.400 ;
  LAYER metal1 ;
  RECT 463.540 763.280 467.080 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 454.860 763.280 458.400 764.400 ;
  LAYER metal3 ;
  RECT 454.860 763.280 458.400 764.400 ;
  LAYER metal2 ;
  RECT 454.860 763.280 458.400 764.400 ;
  LAYER metal1 ;
  RECT 454.860 763.280 458.400 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 446.180 763.280 449.720 764.400 ;
  LAYER metal3 ;
  RECT 446.180 763.280 449.720 764.400 ;
  LAYER metal2 ;
  RECT 446.180 763.280 449.720 764.400 ;
  LAYER metal1 ;
  RECT 446.180 763.280 449.720 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 402.780 763.280 406.320 764.400 ;
  LAYER metal3 ;
  RECT 402.780 763.280 406.320 764.400 ;
  LAYER metal2 ;
  RECT 402.780 763.280 406.320 764.400 ;
  LAYER metal1 ;
  RECT 402.780 763.280 406.320 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 394.100 763.280 397.640 764.400 ;
  LAYER metal3 ;
  RECT 394.100 763.280 397.640 764.400 ;
  LAYER metal2 ;
  RECT 394.100 763.280 397.640 764.400 ;
  LAYER metal1 ;
  RECT 394.100 763.280 397.640 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 385.420 763.280 388.960 764.400 ;
  LAYER metal3 ;
  RECT 385.420 763.280 388.960 764.400 ;
  LAYER metal2 ;
  RECT 385.420 763.280 388.960 764.400 ;
  LAYER metal1 ;
  RECT 385.420 763.280 388.960 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 376.740 763.280 380.280 764.400 ;
  LAYER metal3 ;
  RECT 376.740 763.280 380.280 764.400 ;
  LAYER metal2 ;
  RECT 376.740 763.280 380.280 764.400 ;
  LAYER metal1 ;
  RECT 376.740 763.280 380.280 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 368.060 763.280 371.600 764.400 ;
  LAYER metal3 ;
  RECT 368.060 763.280 371.600 764.400 ;
  LAYER metal2 ;
  RECT 368.060 763.280 371.600 764.400 ;
  LAYER metal1 ;
  RECT 368.060 763.280 371.600 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 359.380 763.280 362.920 764.400 ;
  LAYER metal3 ;
  RECT 359.380 763.280 362.920 764.400 ;
  LAYER metal2 ;
  RECT 359.380 763.280 362.920 764.400 ;
  LAYER metal1 ;
  RECT 359.380 763.280 362.920 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.980 763.280 319.520 764.400 ;
  LAYER metal3 ;
  RECT 315.980 763.280 319.520 764.400 ;
  LAYER metal2 ;
  RECT 315.980 763.280 319.520 764.400 ;
  LAYER metal1 ;
  RECT 315.980 763.280 319.520 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 307.300 763.280 310.840 764.400 ;
  LAYER metal3 ;
  RECT 307.300 763.280 310.840 764.400 ;
  LAYER metal2 ;
  RECT 307.300 763.280 310.840 764.400 ;
  LAYER metal1 ;
  RECT 307.300 763.280 310.840 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 298.620 763.280 302.160 764.400 ;
  LAYER metal3 ;
  RECT 298.620 763.280 302.160 764.400 ;
  LAYER metal2 ;
  RECT 298.620 763.280 302.160 764.400 ;
  LAYER metal1 ;
  RECT 298.620 763.280 302.160 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 289.940 763.280 293.480 764.400 ;
  LAYER metal3 ;
  RECT 289.940 763.280 293.480 764.400 ;
  LAYER metal2 ;
  RECT 289.940 763.280 293.480 764.400 ;
  LAYER metal1 ;
  RECT 289.940 763.280 293.480 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 281.260 763.280 284.800 764.400 ;
  LAYER metal3 ;
  RECT 281.260 763.280 284.800 764.400 ;
  LAYER metal2 ;
  RECT 281.260 763.280 284.800 764.400 ;
  LAYER metal1 ;
  RECT 281.260 763.280 284.800 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 272.580 763.280 276.120 764.400 ;
  LAYER metal3 ;
  RECT 272.580 763.280 276.120 764.400 ;
  LAYER metal2 ;
  RECT 272.580 763.280 276.120 764.400 ;
  LAYER metal1 ;
  RECT 272.580 763.280 276.120 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.180 763.280 232.720 764.400 ;
  LAYER metal3 ;
  RECT 229.180 763.280 232.720 764.400 ;
  LAYER metal2 ;
  RECT 229.180 763.280 232.720 764.400 ;
  LAYER metal1 ;
  RECT 229.180 763.280 232.720 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 220.500 763.280 224.040 764.400 ;
  LAYER metal3 ;
  RECT 220.500 763.280 224.040 764.400 ;
  LAYER metal2 ;
  RECT 220.500 763.280 224.040 764.400 ;
  LAYER metal1 ;
  RECT 220.500 763.280 224.040 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 211.820 763.280 215.360 764.400 ;
  LAYER metal3 ;
  RECT 211.820 763.280 215.360 764.400 ;
  LAYER metal2 ;
  RECT 211.820 763.280 215.360 764.400 ;
  LAYER metal1 ;
  RECT 211.820 763.280 215.360 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 203.140 763.280 206.680 764.400 ;
  LAYER metal3 ;
  RECT 203.140 763.280 206.680 764.400 ;
  LAYER metal2 ;
  RECT 203.140 763.280 206.680 764.400 ;
  LAYER metal1 ;
  RECT 203.140 763.280 206.680 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 194.460 763.280 198.000 764.400 ;
  LAYER metal3 ;
  RECT 194.460 763.280 198.000 764.400 ;
  LAYER metal2 ;
  RECT 194.460 763.280 198.000 764.400 ;
  LAYER metal1 ;
  RECT 194.460 763.280 198.000 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 185.780 763.280 189.320 764.400 ;
  LAYER metal3 ;
  RECT 185.780 763.280 189.320 764.400 ;
  LAYER metal2 ;
  RECT 185.780 763.280 189.320 764.400 ;
  LAYER metal1 ;
  RECT 185.780 763.280 189.320 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 142.380 763.280 145.920 764.400 ;
  LAYER metal3 ;
  RECT 142.380 763.280 145.920 764.400 ;
  LAYER metal2 ;
  RECT 142.380 763.280 145.920 764.400 ;
  LAYER metal1 ;
  RECT 142.380 763.280 145.920 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 133.700 763.280 137.240 764.400 ;
  LAYER metal3 ;
  RECT 133.700 763.280 137.240 764.400 ;
  LAYER metal2 ;
  RECT 133.700 763.280 137.240 764.400 ;
  LAYER metal1 ;
  RECT 133.700 763.280 137.240 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 125.020 763.280 128.560 764.400 ;
  LAYER metal3 ;
  RECT 125.020 763.280 128.560 764.400 ;
  LAYER metal2 ;
  RECT 125.020 763.280 128.560 764.400 ;
  LAYER metal1 ;
  RECT 125.020 763.280 128.560 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 116.340 763.280 119.880 764.400 ;
  LAYER metal3 ;
  RECT 116.340 763.280 119.880 764.400 ;
  LAYER metal2 ;
  RECT 116.340 763.280 119.880 764.400 ;
  LAYER metal1 ;
  RECT 116.340 763.280 119.880 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 107.660 763.280 111.200 764.400 ;
  LAYER metal3 ;
  RECT 107.660 763.280 111.200 764.400 ;
  LAYER metal2 ;
  RECT 107.660 763.280 111.200 764.400 ;
  LAYER metal1 ;
  RECT 107.660 763.280 111.200 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 98.980 763.280 102.520 764.400 ;
  LAYER metal3 ;
  RECT 98.980 763.280 102.520 764.400 ;
  LAYER metal2 ;
  RECT 98.980 763.280 102.520 764.400 ;
  LAYER metal1 ;
  RECT 98.980 763.280 102.520 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 55.580 763.280 59.120 764.400 ;
  LAYER metal3 ;
  RECT 55.580 763.280 59.120 764.400 ;
  LAYER metal2 ;
  RECT 55.580 763.280 59.120 764.400 ;
  LAYER metal1 ;
  RECT 55.580 763.280 59.120 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 46.900 763.280 50.440 764.400 ;
  LAYER metal3 ;
  RECT 46.900 763.280 50.440 764.400 ;
  LAYER metal2 ;
  RECT 46.900 763.280 50.440 764.400 ;
  LAYER metal1 ;
  RECT 46.900 763.280 50.440 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 38.220 763.280 41.760 764.400 ;
  LAYER metal3 ;
  RECT 38.220 763.280 41.760 764.400 ;
  LAYER metal2 ;
  RECT 38.220 763.280 41.760 764.400 ;
  LAYER metal1 ;
  RECT 38.220 763.280 41.760 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 29.540 763.280 33.080 764.400 ;
  LAYER metal3 ;
  RECT 29.540 763.280 33.080 764.400 ;
  LAYER metal2 ;
  RECT 29.540 763.280 33.080 764.400 ;
  LAYER metal1 ;
  RECT 29.540 763.280 33.080 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 20.860 763.280 24.400 764.400 ;
  LAYER metal3 ;
  RECT 20.860 763.280 24.400 764.400 ;
  LAYER metal2 ;
  RECT 20.860 763.280 24.400 764.400 ;
  LAYER metal1 ;
  RECT 20.860 763.280 24.400 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.180 763.280 15.720 764.400 ;
  LAYER metal3 ;
  RECT 12.180 763.280 15.720 764.400 ;
  LAYER metal2 ;
  RECT 12.180 763.280 15.720 764.400 ;
  LAYER metal1 ;
  RECT 12.180 763.280 15.720 764.400 ;
 END
 PORT
  LAYER metal4 ;
  RECT 965.120 0.000 968.660 1.120 ;
  LAYER metal3 ;
  RECT 965.120 0.000 968.660 1.120 ;
  LAYER metal2 ;
  RECT 965.120 0.000 968.660 1.120 ;
  LAYER metal1 ;
  RECT 965.120 0.000 968.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 956.440 0.000 959.980 1.120 ;
  LAYER metal3 ;
  RECT 956.440 0.000 959.980 1.120 ;
  LAYER metal2 ;
  RECT 956.440 0.000 959.980 1.120 ;
  LAYER metal1 ;
  RECT 956.440 0.000 959.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 947.760 0.000 951.300 1.120 ;
  LAYER metal3 ;
  RECT 947.760 0.000 951.300 1.120 ;
  LAYER metal2 ;
  RECT 947.760 0.000 951.300 1.120 ;
  LAYER metal1 ;
  RECT 947.760 0.000 951.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 939.080 0.000 942.620 1.120 ;
  LAYER metal3 ;
  RECT 939.080 0.000 942.620 1.120 ;
  LAYER metal2 ;
  RECT 939.080 0.000 942.620 1.120 ;
  LAYER metal1 ;
  RECT 939.080 0.000 942.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 930.400 0.000 933.940 1.120 ;
  LAYER metal3 ;
  RECT 930.400 0.000 933.940 1.120 ;
  LAYER metal2 ;
  RECT 930.400 0.000 933.940 1.120 ;
  LAYER metal1 ;
  RECT 930.400 0.000 933.940 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 921.720 0.000 925.260 1.120 ;
  LAYER metal3 ;
  RECT 921.720 0.000 925.260 1.120 ;
  LAYER metal2 ;
  RECT 921.720 0.000 925.260 1.120 ;
  LAYER metal1 ;
  RECT 921.720 0.000 925.260 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 878.320 0.000 881.860 1.120 ;
  LAYER metal3 ;
  RECT 878.320 0.000 881.860 1.120 ;
  LAYER metal2 ;
  RECT 878.320 0.000 881.860 1.120 ;
  LAYER metal1 ;
  RECT 878.320 0.000 881.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 869.640 0.000 873.180 1.120 ;
  LAYER metal3 ;
  RECT 869.640 0.000 873.180 1.120 ;
  LAYER metal2 ;
  RECT 869.640 0.000 873.180 1.120 ;
  LAYER metal1 ;
  RECT 869.640 0.000 873.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 860.960 0.000 864.500 1.120 ;
  LAYER metal3 ;
  RECT 860.960 0.000 864.500 1.120 ;
  LAYER metal2 ;
  RECT 860.960 0.000 864.500 1.120 ;
  LAYER metal1 ;
  RECT 860.960 0.000 864.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal3 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal2 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal1 ;
  RECT 852.280 0.000 855.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 843.600 0.000 847.140 1.120 ;
  LAYER metal3 ;
  RECT 843.600 0.000 847.140 1.120 ;
  LAYER metal2 ;
  RECT 843.600 0.000 847.140 1.120 ;
  LAYER metal1 ;
  RECT 843.600 0.000 847.140 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal3 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal2 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal1 ;
  RECT 834.920 0.000 838.460 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 774.160 0.000 777.700 1.120 ;
  LAYER metal3 ;
  RECT 774.160 0.000 777.700 1.120 ;
  LAYER metal2 ;
  RECT 774.160 0.000 777.700 1.120 ;
  LAYER metal1 ;
  RECT 774.160 0.000 777.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 765.480 0.000 769.020 1.120 ;
  LAYER metal3 ;
  RECT 765.480 0.000 769.020 1.120 ;
  LAYER metal2 ;
  RECT 765.480 0.000 769.020 1.120 ;
  LAYER metal1 ;
  RECT 765.480 0.000 769.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 756.800 0.000 760.340 1.120 ;
  LAYER metal3 ;
  RECT 756.800 0.000 760.340 1.120 ;
  LAYER metal2 ;
  RECT 756.800 0.000 760.340 1.120 ;
  LAYER metal1 ;
  RECT 756.800 0.000 760.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 748.120 0.000 751.660 1.120 ;
  LAYER metal3 ;
  RECT 748.120 0.000 751.660 1.120 ;
  LAYER metal2 ;
  RECT 748.120 0.000 751.660 1.120 ;
  LAYER metal1 ;
  RECT 748.120 0.000 751.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 739.440 0.000 742.980 1.120 ;
  LAYER metal3 ;
  RECT 739.440 0.000 742.980 1.120 ;
  LAYER metal2 ;
  RECT 739.440 0.000 742.980 1.120 ;
  LAYER metal1 ;
  RECT 739.440 0.000 742.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 730.760 0.000 734.300 1.120 ;
  LAYER metal3 ;
  RECT 730.760 0.000 734.300 1.120 ;
  LAYER metal2 ;
  RECT 730.760 0.000 734.300 1.120 ;
  LAYER metal1 ;
  RECT 730.760 0.000 734.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 687.360 0.000 690.900 1.120 ;
  LAYER metal3 ;
  RECT 687.360 0.000 690.900 1.120 ;
  LAYER metal2 ;
  RECT 687.360 0.000 690.900 1.120 ;
  LAYER metal1 ;
  RECT 687.360 0.000 690.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER metal3 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER metal2 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER metal1 ;
  RECT 678.680 0.000 682.220 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 670.000 0.000 673.540 1.120 ;
  LAYER metal3 ;
  RECT 670.000 0.000 673.540 1.120 ;
  LAYER metal2 ;
  RECT 670.000 0.000 673.540 1.120 ;
  LAYER metal1 ;
  RECT 670.000 0.000 673.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 661.320 0.000 664.860 1.120 ;
  LAYER metal3 ;
  RECT 661.320 0.000 664.860 1.120 ;
  LAYER metal2 ;
  RECT 661.320 0.000 664.860 1.120 ;
  LAYER metal1 ;
  RECT 661.320 0.000 664.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 652.640 0.000 656.180 1.120 ;
  LAYER metal3 ;
  RECT 652.640 0.000 656.180 1.120 ;
  LAYER metal2 ;
  RECT 652.640 0.000 656.180 1.120 ;
  LAYER metal1 ;
  RECT 652.640 0.000 656.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 643.960 0.000 647.500 1.120 ;
  LAYER metal3 ;
  RECT 643.960 0.000 647.500 1.120 ;
  LAYER metal2 ;
  RECT 643.960 0.000 647.500 1.120 ;
  LAYER metal1 ;
  RECT 643.960 0.000 647.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 600.560 0.000 604.100 1.120 ;
  LAYER metal3 ;
  RECT 600.560 0.000 604.100 1.120 ;
  LAYER metal2 ;
  RECT 600.560 0.000 604.100 1.120 ;
  LAYER metal1 ;
  RECT 600.560 0.000 604.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER metal3 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER metal2 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER metal1 ;
  RECT 591.880 0.000 595.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 583.200 0.000 586.740 1.120 ;
  LAYER metal3 ;
  RECT 583.200 0.000 586.740 1.120 ;
  LAYER metal2 ;
  RECT 583.200 0.000 586.740 1.120 ;
  LAYER metal1 ;
  RECT 583.200 0.000 586.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal3 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal2 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal1 ;
  RECT 570.180 0.000 573.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 534.220 0.000 537.760 1.120 ;
  LAYER metal3 ;
  RECT 534.220 0.000 537.760 1.120 ;
  LAYER metal2 ;
  RECT 534.220 0.000 537.760 1.120 ;
  LAYER metal1 ;
  RECT 534.220 0.000 537.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 503.840 0.000 507.380 1.120 ;
  LAYER metal3 ;
  RECT 503.840 0.000 507.380 1.120 ;
  LAYER metal2 ;
  RECT 503.840 0.000 507.380 1.120 ;
  LAYER metal1 ;
  RECT 503.840 0.000 507.380 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 439.360 0.000 442.900 1.120 ;
  LAYER metal3 ;
  RECT 439.360 0.000 442.900 1.120 ;
  LAYER metal2 ;
  RECT 439.360 0.000 442.900 1.120 ;
  LAYER metal1 ;
  RECT 439.360 0.000 442.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 430.680 0.000 434.220 1.120 ;
  LAYER metal3 ;
  RECT 430.680 0.000 434.220 1.120 ;
  LAYER metal2 ;
  RECT 430.680 0.000 434.220 1.120 ;
  LAYER metal1 ;
  RECT 430.680 0.000 434.220 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 422.000 0.000 425.540 1.120 ;
  LAYER metal3 ;
  RECT 422.000 0.000 425.540 1.120 ;
  LAYER metal2 ;
  RECT 422.000 0.000 425.540 1.120 ;
  LAYER metal1 ;
  RECT 422.000 0.000 425.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 413.320 0.000 416.860 1.120 ;
  LAYER metal3 ;
  RECT 413.320 0.000 416.860 1.120 ;
  LAYER metal2 ;
  RECT 413.320 0.000 416.860 1.120 ;
  LAYER metal1 ;
  RECT 413.320 0.000 416.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 404.640 0.000 408.180 1.120 ;
  LAYER metal3 ;
  RECT 404.640 0.000 408.180 1.120 ;
  LAYER metal2 ;
  RECT 404.640 0.000 408.180 1.120 ;
  LAYER metal1 ;
  RECT 404.640 0.000 408.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 395.960 0.000 399.500 1.120 ;
  LAYER metal3 ;
  RECT 395.960 0.000 399.500 1.120 ;
  LAYER metal2 ;
  RECT 395.960 0.000 399.500 1.120 ;
  LAYER metal1 ;
  RECT 395.960 0.000 399.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 352.560 0.000 356.100 1.120 ;
  LAYER metal3 ;
  RECT 352.560 0.000 356.100 1.120 ;
  LAYER metal2 ;
  RECT 352.560 0.000 356.100 1.120 ;
  LAYER metal1 ;
  RECT 352.560 0.000 356.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 343.880 0.000 347.420 1.120 ;
  LAYER metal3 ;
  RECT 343.880 0.000 347.420 1.120 ;
  LAYER metal2 ;
  RECT 343.880 0.000 347.420 1.120 ;
  LAYER metal1 ;
  RECT 343.880 0.000 347.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 335.200 0.000 338.740 1.120 ;
  LAYER metal3 ;
  RECT 335.200 0.000 338.740 1.120 ;
  LAYER metal2 ;
  RECT 335.200 0.000 338.740 1.120 ;
  LAYER metal1 ;
  RECT 335.200 0.000 338.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal3 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal2 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal1 ;
  RECT 326.520 0.000 330.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 317.840 0.000 321.380 1.120 ;
  LAYER metal3 ;
  RECT 317.840 0.000 321.380 1.120 ;
  LAYER metal2 ;
  RECT 317.840 0.000 321.380 1.120 ;
  LAYER metal1 ;
  RECT 317.840 0.000 321.380 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 309.160 0.000 312.700 1.120 ;
  LAYER metal3 ;
  RECT 309.160 0.000 312.700 1.120 ;
  LAYER metal2 ;
  RECT 309.160 0.000 312.700 1.120 ;
  LAYER metal1 ;
  RECT 309.160 0.000 312.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 265.760 0.000 269.300 1.120 ;
  LAYER metal3 ;
  RECT 265.760 0.000 269.300 1.120 ;
  LAYER metal2 ;
  RECT 265.760 0.000 269.300 1.120 ;
  LAYER metal1 ;
  RECT 265.760 0.000 269.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal3 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal2 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal1 ;
  RECT 253.360 0.000 256.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 231.040 0.000 234.580 1.120 ;
  LAYER metal3 ;
  RECT 231.040 0.000 234.580 1.120 ;
  LAYER metal2 ;
  RECT 231.040 0.000 234.580 1.120 ;
  LAYER metal1 ;
  RECT 231.040 0.000 234.580 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 222.360 0.000 225.900 1.120 ;
  LAYER metal3 ;
  RECT 222.360 0.000 225.900 1.120 ;
  LAYER metal2 ;
  RECT 222.360 0.000 225.900 1.120 ;
  LAYER metal1 ;
  RECT 222.360 0.000 225.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 213.680 0.000 217.220 1.120 ;
  LAYER metal3 ;
  RECT 213.680 0.000 217.220 1.120 ;
  LAYER metal2 ;
  RECT 213.680 0.000 217.220 1.120 ;
  LAYER metal1 ;
  RECT 213.680 0.000 217.220 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 205.000 0.000 208.540 1.120 ;
  LAYER metal3 ;
  RECT 205.000 0.000 208.540 1.120 ;
  LAYER metal2 ;
  RECT 205.000 0.000 208.540 1.120 ;
  LAYER metal1 ;
  RECT 205.000 0.000 208.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 161.600 0.000 165.140 1.120 ;
  LAYER metal3 ;
  RECT 161.600 0.000 165.140 1.120 ;
  LAYER metal2 ;
  RECT 161.600 0.000 165.140 1.120 ;
  LAYER metal1 ;
  RECT 161.600 0.000 165.140 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 152.920 0.000 156.460 1.120 ;
  LAYER metal3 ;
  RECT 152.920 0.000 156.460 1.120 ;
  LAYER metal2 ;
  RECT 152.920 0.000 156.460 1.120 ;
  LAYER metal1 ;
  RECT 152.920 0.000 156.460 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 144.240 0.000 147.780 1.120 ;
  LAYER metal3 ;
  RECT 144.240 0.000 147.780 1.120 ;
  LAYER metal2 ;
  RECT 144.240 0.000 147.780 1.120 ;
  LAYER metal1 ;
  RECT 144.240 0.000 147.780 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 135.560 0.000 139.100 1.120 ;
  LAYER metal3 ;
  RECT 135.560 0.000 139.100 1.120 ;
  LAYER metal2 ;
  RECT 135.560 0.000 139.100 1.120 ;
  LAYER metal1 ;
  RECT 135.560 0.000 139.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 118.200 0.000 121.740 1.120 ;
  LAYER metal3 ;
  RECT 118.200 0.000 121.740 1.120 ;
  LAYER metal2 ;
  RECT 118.200 0.000 121.740 1.120 ;
  LAYER metal1 ;
  RECT 118.200 0.000 121.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 74.800 0.000 78.340 1.120 ;
  LAYER metal3 ;
  RECT 74.800 0.000 78.340 1.120 ;
  LAYER metal2 ;
  RECT 74.800 0.000 78.340 1.120 ;
  LAYER metal1 ;
  RECT 74.800 0.000 78.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 66.120 0.000 69.660 1.120 ;
  LAYER metal3 ;
  RECT 66.120 0.000 69.660 1.120 ;
  LAYER metal2 ;
  RECT 66.120 0.000 69.660 1.120 ;
  LAYER metal1 ;
  RECT 66.120 0.000 69.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER metal3 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER metal2 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER metal1 ;
  RECT 57.440 0.000 60.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER metal3 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER metal2 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER metal1 ;
  RECT 48.760 0.000 52.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER metal3 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER metal2 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER metal1 ;
  RECT 40.080 0.000 43.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.228 ;
 PORT
  LAYER metal4 ;
  RECT 802.340 0.000 803.460 1.120 ;
  LAYER metal3 ;
  RECT 802.340 0.000 803.460 1.120 ;
  LAYER metal2 ;
  RECT 802.340 0.000 803.460 1.120 ;
  LAYER metal1 ;
  RECT 802.340 0.000 803.460 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.079 ;
 PORT
  LAYER metal4 ;
  RECT 794.280 0.000 795.400 1.120 ;
  LAYER metal3 ;
  RECT 794.280 0.000 795.400 1.120 ;
  LAYER metal2 ;
  RECT 794.280 0.000 795.400 1.120 ;
  LAYER metal1 ;
  RECT 794.280 0.000 795.400 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.228 ;
 PORT
  LAYER metal4 ;
  RECT 789.320 0.000 790.440 1.120 ;
  LAYER metal3 ;
  RECT 789.320 0.000 790.440 1.120 ;
  LAYER metal2 ;
  RECT 789.320 0.000 790.440 1.120 ;
  LAYER metal1 ;
  RECT 789.320 0.000 790.440 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.079 ;
 PORT
  LAYER metal4 ;
  RECT 781.260 0.000 782.380 1.120 ;
  LAYER metal3 ;
  RECT 781.260 0.000 782.380 1.120 ;
  LAYER metal2 ;
  RECT 781.260 0.000 782.380 1.120 ;
  LAYER metal1 ;
  RECT 781.260 0.000 782.380 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.228 ;
 PORT
  LAYER metal4 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER metal3 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER metal2 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER metal1 ;
  RECT 576.660 0.000 577.780 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.079 ;
 PORT
  LAYER metal4 ;
  RECT 567.980 0.000 569.100 1.120 ;
  LAYER metal3 ;
  RECT 567.980 0.000 569.100 1.120 ;
  LAYER metal2 ;
  RECT 567.980 0.000 569.100 1.120 ;
  LAYER metal1 ;
  RECT 567.980 0.000 569.100 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.228 ;
 PORT
  LAYER metal4 ;
  RECT 563.020 0.000 564.140 1.120 ;
  LAYER metal3 ;
  RECT 563.020 0.000 564.140 1.120 ;
  LAYER metal2 ;
  RECT 563.020 0.000 564.140 1.120 ;
  LAYER metal1 ;
  RECT 563.020 0.000 564.140 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.079 ;
 PORT
  LAYER metal4 ;
  RECT 554.960 0.000 556.080 1.120 ;
  LAYER metal3 ;
  RECT 554.960 0.000 556.080 1.120 ;
  LAYER metal2 ;
  RECT 554.960 0.000 556.080 1.120 ;
  LAYER metal1 ;
  RECT 554.960 0.000 556.080 1.120 ;
 END
END DI4
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 549.380 0.000 550.500 1.120 ;
  LAYER metal3 ;
  RECT 549.380 0.000 550.500 1.120 ;
  LAYER metal2 ;
  RECT 549.380 0.000 550.500 1.120 ;
  LAYER metal1 ;
  RECT 549.380 0.000 550.500 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 547.520 0.000 548.640 1.120 ;
  LAYER metal3 ;
  RECT 547.520 0.000 548.640 1.120 ;
  LAYER metal2 ;
  RECT 547.520 0.000 548.640 1.120 ;
  LAYER metal1 ;
  RECT 547.520 0.000 548.640 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER metal4 ;
  RECT 542.560 0.000 543.680 1.120 ;
  LAYER metal3 ;
  RECT 542.560 0.000 543.680 1.120 ;
  LAYER metal2 ;
  RECT 542.560 0.000 543.680 1.120 ;
  LAYER metal1 ;
  RECT 542.560 0.000 543.680 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER metal4 ;
  RECT 540.700 0.000 541.820 1.120 ;
  LAYER metal3 ;
  RECT 540.700 0.000 541.820 1.120 ;
  LAYER metal2 ;
  RECT 540.700 0.000 541.820 1.120 ;
  LAYER metal1 ;
  RECT 540.700 0.000 541.820 1.120 ;
 END
END CS
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 538.840 0.000 539.960 1.120 ;
  LAYER metal3 ;
  RECT 538.840 0.000 539.960 1.120 ;
  LAYER metal2 ;
  RECT 538.840 0.000 539.960 1.120 ;
  LAYER metal1 ;
  RECT 538.840 0.000 539.960 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 532.020 0.000 533.140 1.120 ;
  LAYER metal3 ;
  RECT 532.020 0.000 533.140 1.120 ;
  LAYER metal2 ;
  RECT 532.020 0.000 533.140 1.120 ;
  LAYER metal1 ;
  RECT 532.020 0.000 533.140 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 529.540 0.000 530.660 1.120 ;
  LAYER metal3 ;
  RECT 529.540 0.000 530.660 1.120 ;
  LAYER metal2 ;
  RECT 529.540 0.000 530.660 1.120 ;
  LAYER metal1 ;
  RECT 529.540 0.000 530.660 1.120 ;
 END
END A5
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 519.000 0.000 520.120 1.120 ;
  LAYER metal3 ;
  RECT 519.000 0.000 520.120 1.120 ;
  LAYER metal2 ;
  RECT 519.000 0.000 520.120 1.120 ;
  LAYER metal1 ;
  RECT 519.000 0.000 520.120 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER metal4 ;
  RECT 515.900 0.000 517.020 1.120 ;
  LAYER metal3 ;
  RECT 515.900 0.000 517.020 1.120 ;
  LAYER metal2 ;
  RECT 515.900 0.000 517.020 1.120 ;
  LAYER metal1 ;
  RECT 515.900 0.000 517.020 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 514.040 0.000 515.160 1.120 ;
  LAYER metal3 ;
  RECT 514.040 0.000 515.160 1.120 ;
  LAYER metal2 ;
  RECT 514.040 0.000 515.160 1.120 ;
  LAYER metal1 ;
  RECT 514.040 0.000 515.160 1.120 ;
 END
END A0
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER metal3 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER metal2 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER metal1 ;
  RECT 509.700 0.000 510.820 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 501.640 0.000 502.760 1.120 ;
  LAYER metal3 ;
  RECT 501.640 0.000 502.760 1.120 ;
  LAYER metal2 ;
  RECT 501.640 0.000 502.760 1.120 ;
  LAYER metal1 ;
  RECT 501.640 0.000 502.760 1.120 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 499.160 0.000 500.280 1.120 ;
  LAYER metal3 ;
  RECT 499.160 0.000 500.280 1.120 ;
  LAYER metal2 ;
  RECT 499.160 0.000 500.280 1.120 ;
  LAYER metal1 ;
  RECT 499.160 0.000 500.280 1.120 ;
 END
END A8
PIN A9
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 491.100 0.000 492.220 1.120 ;
  LAYER metal3 ;
  RECT 491.100 0.000 492.220 1.120 ;
  LAYER metal2 ;
  RECT 491.100 0.000 492.220 1.120 ;
  LAYER metal1 ;
  RECT 491.100 0.000 492.220 1.120 ;
 END
END A9
PIN A10
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal3 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal2 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal1 ;
  RECT 488.000 0.000 489.120 1.120 ;
 END
END A10
PIN A11
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 480.560 0.000 481.680 1.120 ;
  LAYER metal3 ;
  RECT 480.560 0.000 481.680 1.120 ;
  LAYER metal2 ;
  RECT 480.560 0.000 481.680 1.120 ;
  LAYER metal1 ;
  RECT 480.560 0.000 481.680 1.120 ;
 END
END A11
PIN A12
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER metal3 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER metal2 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER metal1 ;
  RECT 477.460 0.000 478.580 1.120 ;
 END
END A12
PIN A13
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 470.020 0.000 471.140 1.120 ;
  LAYER metal3 ;
  RECT 470.020 0.000 471.140 1.120 ;
  LAYER metal2 ;
  RECT 470.020 0.000 471.140 1.120 ;
  LAYER metal1 ;
  RECT 470.020 0.000 471.140 1.120 ;
 END
END A13
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.228 ;
 PORT
  LAYER metal4 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal3 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal2 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal1 ;
  RECT 259.220 0.000 260.340 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.079 ;
 PORT
  LAYER metal4 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal3 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal2 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal1 ;
  RECT 251.160 0.000 252.280 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.228 ;
 PORT
  LAYER metal4 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal3 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal2 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal1 ;
  RECT 246.200 0.000 247.320 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.079 ;
 PORT
  LAYER metal4 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal3 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal2 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal1 ;
  RECT 237.520 0.000 238.640 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.228 ;
 PORT
  LAYER metal4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.079 ;
 PORT
  LAYER metal4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.228 ;
 PORT
  LAYER metal4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.079 ;
 PORT
  LAYER metal4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 1015.560 764.400 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 1015.560 764.400 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 1015.560 764.400 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 1015.560 764.400 ;
  LAYER via ;
  RECT 0.000 0.140 1015.560 764.400 ;
  LAYER via2 ;
  RECT 0.000 0.140 1015.560 764.400 ;
  LAYER via3 ;
  RECT 0.000 0.140 1015.560 764.400 ;
END
END Img
END LIBRARY



