# 
#              Synchronous Dual Port SRAM Compiler 
# 
#                    UMC 0.18um Generic Logic Process 
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : SRAM_1296X20
#       Words            : 1296
#       Bits             : 20
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2023/10/20 23:57:47
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SRAM_1296X20
CLASS BLOCK ;
FOREIGN SRAM_1296X20 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 674.560 BY 647.920 ;
SYMMETRY x y r90 ;
SITE core_5040 ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal5 ;
  RECT 673.440 634.820 674.560 638.060 ;
  LAYER metal4 ;
  RECT 673.440 634.820 674.560 638.060 ;
  LAYER metal3 ;
  RECT 673.440 634.820 674.560 638.060 ;
  LAYER metal2 ;
  RECT 673.440 634.820 674.560 638.060 ;
  LAYER metal1 ;
  RECT 673.440 634.820 674.560 638.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 595.620 674.560 598.860 ;
  LAYER metal4 ;
  RECT 673.440 595.620 674.560 598.860 ;
  LAYER metal3 ;
  RECT 673.440 595.620 674.560 598.860 ;
  LAYER metal2 ;
  RECT 673.440 595.620 674.560 598.860 ;
  LAYER metal1 ;
  RECT 673.440 595.620 674.560 598.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 587.780 674.560 591.020 ;
  LAYER metal4 ;
  RECT 673.440 587.780 674.560 591.020 ;
  LAYER metal3 ;
  RECT 673.440 587.780 674.560 591.020 ;
  LAYER metal2 ;
  RECT 673.440 587.780 674.560 591.020 ;
  LAYER metal1 ;
  RECT 673.440 587.780 674.560 591.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 579.940 674.560 583.180 ;
  LAYER metal4 ;
  RECT 673.440 579.940 674.560 583.180 ;
  LAYER metal3 ;
  RECT 673.440 579.940 674.560 583.180 ;
  LAYER metal2 ;
  RECT 673.440 579.940 674.560 583.180 ;
  LAYER metal1 ;
  RECT 673.440 579.940 674.560 583.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 572.100 674.560 575.340 ;
  LAYER metal4 ;
  RECT 673.440 572.100 674.560 575.340 ;
  LAYER metal3 ;
  RECT 673.440 572.100 674.560 575.340 ;
  LAYER metal2 ;
  RECT 673.440 572.100 674.560 575.340 ;
  LAYER metal1 ;
  RECT 673.440 572.100 674.560 575.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 564.260 674.560 567.500 ;
  LAYER metal4 ;
  RECT 673.440 564.260 674.560 567.500 ;
  LAYER metal3 ;
  RECT 673.440 564.260 674.560 567.500 ;
  LAYER metal2 ;
  RECT 673.440 564.260 674.560 567.500 ;
  LAYER metal1 ;
  RECT 673.440 564.260 674.560 567.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 556.420 674.560 559.660 ;
  LAYER metal4 ;
  RECT 673.440 556.420 674.560 559.660 ;
  LAYER metal3 ;
  RECT 673.440 556.420 674.560 559.660 ;
  LAYER metal2 ;
  RECT 673.440 556.420 674.560 559.660 ;
  LAYER metal1 ;
  RECT 673.440 556.420 674.560 559.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 517.220 674.560 520.460 ;
  LAYER metal4 ;
  RECT 673.440 517.220 674.560 520.460 ;
  LAYER metal3 ;
  RECT 673.440 517.220 674.560 520.460 ;
  LAYER metal2 ;
  RECT 673.440 517.220 674.560 520.460 ;
  LAYER metal1 ;
  RECT 673.440 517.220 674.560 520.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 509.380 674.560 512.620 ;
  LAYER metal4 ;
  RECT 673.440 509.380 674.560 512.620 ;
  LAYER metal3 ;
  RECT 673.440 509.380 674.560 512.620 ;
  LAYER metal2 ;
  RECT 673.440 509.380 674.560 512.620 ;
  LAYER metal1 ;
  RECT 673.440 509.380 674.560 512.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 501.540 674.560 504.780 ;
  LAYER metal4 ;
  RECT 673.440 501.540 674.560 504.780 ;
  LAYER metal3 ;
  RECT 673.440 501.540 674.560 504.780 ;
  LAYER metal2 ;
  RECT 673.440 501.540 674.560 504.780 ;
  LAYER metal1 ;
  RECT 673.440 501.540 674.560 504.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 493.700 674.560 496.940 ;
  LAYER metal4 ;
  RECT 673.440 493.700 674.560 496.940 ;
  LAYER metal3 ;
  RECT 673.440 493.700 674.560 496.940 ;
  LAYER metal2 ;
  RECT 673.440 493.700 674.560 496.940 ;
  LAYER metal1 ;
  RECT 673.440 493.700 674.560 496.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 485.860 674.560 489.100 ;
  LAYER metal4 ;
  RECT 673.440 485.860 674.560 489.100 ;
  LAYER metal3 ;
  RECT 673.440 485.860 674.560 489.100 ;
  LAYER metal2 ;
  RECT 673.440 485.860 674.560 489.100 ;
  LAYER metal1 ;
  RECT 673.440 485.860 674.560 489.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 478.020 674.560 481.260 ;
  LAYER metal4 ;
  RECT 673.440 478.020 674.560 481.260 ;
  LAYER metal3 ;
  RECT 673.440 478.020 674.560 481.260 ;
  LAYER metal2 ;
  RECT 673.440 478.020 674.560 481.260 ;
  LAYER metal1 ;
  RECT 673.440 478.020 674.560 481.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 438.820 674.560 442.060 ;
  LAYER metal4 ;
  RECT 673.440 438.820 674.560 442.060 ;
  LAYER metal3 ;
  RECT 673.440 438.820 674.560 442.060 ;
  LAYER metal2 ;
  RECT 673.440 438.820 674.560 442.060 ;
  LAYER metal1 ;
  RECT 673.440 438.820 674.560 442.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 430.980 674.560 434.220 ;
  LAYER metal4 ;
  RECT 673.440 430.980 674.560 434.220 ;
  LAYER metal3 ;
  RECT 673.440 430.980 674.560 434.220 ;
  LAYER metal2 ;
  RECT 673.440 430.980 674.560 434.220 ;
  LAYER metal1 ;
  RECT 673.440 430.980 674.560 434.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 423.140 674.560 426.380 ;
  LAYER metal4 ;
  RECT 673.440 423.140 674.560 426.380 ;
  LAYER metal3 ;
  RECT 673.440 423.140 674.560 426.380 ;
  LAYER metal2 ;
  RECT 673.440 423.140 674.560 426.380 ;
  LAYER metal1 ;
  RECT 673.440 423.140 674.560 426.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 415.300 674.560 418.540 ;
  LAYER metal4 ;
  RECT 673.440 415.300 674.560 418.540 ;
  LAYER metal3 ;
  RECT 673.440 415.300 674.560 418.540 ;
  LAYER metal2 ;
  RECT 673.440 415.300 674.560 418.540 ;
  LAYER metal1 ;
  RECT 673.440 415.300 674.560 418.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 407.460 674.560 410.700 ;
  LAYER metal4 ;
  RECT 673.440 407.460 674.560 410.700 ;
  LAYER metal3 ;
  RECT 673.440 407.460 674.560 410.700 ;
  LAYER metal2 ;
  RECT 673.440 407.460 674.560 410.700 ;
  LAYER metal1 ;
  RECT 673.440 407.460 674.560 410.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 399.620 674.560 402.860 ;
  LAYER metal4 ;
  RECT 673.440 399.620 674.560 402.860 ;
  LAYER metal3 ;
  RECT 673.440 399.620 674.560 402.860 ;
  LAYER metal2 ;
  RECT 673.440 399.620 674.560 402.860 ;
  LAYER metal1 ;
  RECT 673.440 399.620 674.560 402.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 360.420 674.560 363.660 ;
  LAYER metal4 ;
  RECT 673.440 360.420 674.560 363.660 ;
  LAYER metal3 ;
  RECT 673.440 360.420 674.560 363.660 ;
  LAYER metal2 ;
  RECT 673.440 360.420 674.560 363.660 ;
  LAYER metal1 ;
  RECT 673.440 360.420 674.560 363.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 352.580 674.560 355.820 ;
  LAYER metal4 ;
  RECT 673.440 352.580 674.560 355.820 ;
  LAYER metal3 ;
  RECT 673.440 352.580 674.560 355.820 ;
  LAYER metal2 ;
  RECT 673.440 352.580 674.560 355.820 ;
  LAYER metal1 ;
  RECT 673.440 352.580 674.560 355.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 344.740 674.560 347.980 ;
  LAYER metal4 ;
  RECT 673.440 344.740 674.560 347.980 ;
  LAYER metal3 ;
  RECT 673.440 344.740 674.560 347.980 ;
  LAYER metal2 ;
  RECT 673.440 344.740 674.560 347.980 ;
  LAYER metal1 ;
  RECT 673.440 344.740 674.560 347.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 336.900 674.560 340.140 ;
  LAYER metal4 ;
  RECT 673.440 336.900 674.560 340.140 ;
  LAYER metal3 ;
  RECT 673.440 336.900 674.560 340.140 ;
  LAYER metal2 ;
  RECT 673.440 336.900 674.560 340.140 ;
  LAYER metal1 ;
  RECT 673.440 336.900 674.560 340.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 329.060 674.560 332.300 ;
  LAYER metal4 ;
  RECT 673.440 329.060 674.560 332.300 ;
  LAYER metal3 ;
  RECT 673.440 329.060 674.560 332.300 ;
  LAYER metal2 ;
  RECT 673.440 329.060 674.560 332.300 ;
  LAYER metal1 ;
  RECT 673.440 329.060 674.560 332.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 321.220 674.560 324.460 ;
  LAYER metal4 ;
  RECT 673.440 321.220 674.560 324.460 ;
  LAYER metal3 ;
  RECT 673.440 321.220 674.560 324.460 ;
  LAYER metal2 ;
  RECT 673.440 321.220 674.560 324.460 ;
  LAYER metal1 ;
  RECT 673.440 321.220 674.560 324.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 282.020 674.560 285.260 ;
  LAYER metal4 ;
  RECT 673.440 282.020 674.560 285.260 ;
  LAYER metal3 ;
  RECT 673.440 282.020 674.560 285.260 ;
  LAYER metal2 ;
  RECT 673.440 282.020 674.560 285.260 ;
  LAYER metal1 ;
  RECT 673.440 282.020 674.560 285.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 274.180 674.560 277.420 ;
  LAYER metal4 ;
  RECT 673.440 274.180 674.560 277.420 ;
  LAYER metal3 ;
  RECT 673.440 274.180 674.560 277.420 ;
  LAYER metal2 ;
  RECT 673.440 274.180 674.560 277.420 ;
  LAYER metal1 ;
  RECT 673.440 274.180 674.560 277.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 266.340 674.560 269.580 ;
  LAYER metal4 ;
  RECT 673.440 266.340 674.560 269.580 ;
  LAYER metal3 ;
  RECT 673.440 266.340 674.560 269.580 ;
  LAYER metal2 ;
  RECT 673.440 266.340 674.560 269.580 ;
  LAYER metal1 ;
  RECT 673.440 266.340 674.560 269.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 258.500 674.560 261.740 ;
  LAYER metal4 ;
  RECT 673.440 258.500 674.560 261.740 ;
  LAYER metal3 ;
  RECT 673.440 258.500 674.560 261.740 ;
  LAYER metal2 ;
  RECT 673.440 258.500 674.560 261.740 ;
  LAYER metal1 ;
  RECT 673.440 258.500 674.560 261.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 250.660 674.560 253.900 ;
  LAYER metal4 ;
  RECT 673.440 250.660 674.560 253.900 ;
  LAYER metal3 ;
  RECT 673.440 250.660 674.560 253.900 ;
  LAYER metal2 ;
  RECT 673.440 250.660 674.560 253.900 ;
  LAYER metal1 ;
  RECT 673.440 250.660 674.560 253.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 242.820 674.560 246.060 ;
  LAYER metal4 ;
  RECT 673.440 242.820 674.560 246.060 ;
  LAYER metal3 ;
  RECT 673.440 242.820 674.560 246.060 ;
  LAYER metal2 ;
  RECT 673.440 242.820 674.560 246.060 ;
  LAYER metal1 ;
  RECT 673.440 242.820 674.560 246.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 203.620 674.560 206.860 ;
  LAYER metal4 ;
  RECT 673.440 203.620 674.560 206.860 ;
  LAYER metal3 ;
  RECT 673.440 203.620 674.560 206.860 ;
  LAYER metal2 ;
  RECT 673.440 203.620 674.560 206.860 ;
  LAYER metal1 ;
  RECT 673.440 203.620 674.560 206.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 195.780 674.560 199.020 ;
  LAYER metal4 ;
  RECT 673.440 195.780 674.560 199.020 ;
  LAYER metal3 ;
  RECT 673.440 195.780 674.560 199.020 ;
  LAYER metal2 ;
  RECT 673.440 195.780 674.560 199.020 ;
  LAYER metal1 ;
  RECT 673.440 195.780 674.560 199.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 187.940 674.560 191.180 ;
  LAYER metal4 ;
  RECT 673.440 187.940 674.560 191.180 ;
  LAYER metal3 ;
  RECT 673.440 187.940 674.560 191.180 ;
  LAYER metal2 ;
  RECT 673.440 187.940 674.560 191.180 ;
  LAYER metal1 ;
  RECT 673.440 187.940 674.560 191.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 180.100 674.560 183.340 ;
  LAYER metal4 ;
  RECT 673.440 180.100 674.560 183.340 ;
  LAYER metal3 ;
  RECT 673.440 180.100 674.560 183.340 ;
  LAYER metal2 ;
  RECT 673.440 180.100 674.560 183.340 ;
  LAYER metal1 ;
  RECT 673.440 180.100 674.560 183.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 172.260 674.560 175.500 ;
  LAYER metal4 ;
  RECT 673.440 172.260 674.560 175.500 ;
  LAYER metal3 ;
  RECT 673.440 172.260 674.560 175.500 ;
  LAYER metal2 ;
  RECT 673.440 172.260 674.560 175.500 ;
  LAYER metal1 ;
  RECT 673.440 172.260 674.560 175.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 164.420 674.560 167.660 ;
  LAYER metal4 ;
  RECT 673.440 164.420 674.560 167.660 ;
  LAYER metal3 ;
  RECT 673.440 164.420 674.560 167.660 ;
  LAYER metal2 ;
  RECT 673.440 164.420 674.560 167.660 ;
  LAYER metal1 ;
  RECT 673.440 164.420 674.560 167.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 125.220 674.560 128.460 ;
  LAYER metal4 ;
  RECT 673.440 125.220 674.560 128.460 ;
  LAYER metal3 ;
  RECT 673.440 125.220 674.560 128.460 ;
  LAYER metal2 ;
  RECT 673.440 125.220 674.560 128.460 ;
  LAYER metal1 ;
  RECT 673.440 125.220 674.560 128.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 117.380 674.560 120.620 ;
  LAYER metal4 ;
  RECT 673.440 117.380 674.560 120.620 ;
  LAYER metal3 ;
  RECT 673.440 117.380 674.560 120.620 ;
  LAYER metal2 ;
  RECT 673.440 117.380 674.560 120.620 ;
  LAYER metal1 ;
  RECT 673.440 117.380 674.560 120.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 109.540 674.560 112.780 ;
  LAYER metal4 ;
  RECT 673.440 109.540 674.560 112.780 ;
  LAYER metal3 ;
  RECT 673.440 109.540 674.560 112.780 ;
  LAYER metal2 ;
  RECT 673.440 109.540 674.560 112.780 ;
  LAYER metal1 ;
  RECT 673.440 109.540 674.560 112.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 101.700 674.560 104.940 ;
  LAYER metal4 ;
  RECT 673.440 101.700 674.560 104.940 ;
  LAYER metal3 ;
  RECT 673.440 101.700 674.560 104.940 ;
  LAYER metal2 ;
  RECT 673.440 101.700 674.560 104.940 ;
  LAYER metal1 ;
  RECT 673.440 101.700 674.560 104.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 93.860 674.560 97.100 ;
  LAYER metal4 ;
  RECT 673.440 93.860 674.560 97.100 ;
  LAYER metal3 ;
  RECT 673.440 93.860 674.560 97.100 ;
  LAYER metal2 ;
  RECT 673.440 93.860 674.560 97.100 ;
  LAYER metal1 ;
  RECT 673.440 93.860 674.560 97.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 86.020 674.560 89.260 ;
  LAYER metal4 ;
  RECT 673.440 86.020 674.560 89.260 ;
  LAYER metal3 ;
  RECT 673.440 86.020 674.560 89.260 ;
  LAYER metal2 ;
  RECT 673.440 86.020 674.560 89.260 ;
  LAYER metal1 ;
  RECT 673.440 86.020 674.560 89.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 46.820 674.560 50.060 ;
  LAYER metal4 ;
  RECT 673.440 46.820 674.560 50.060 ;
  LAYER metal3 ;
  RECT 673.440 46.820 674.560 50.060 ;
  LAYER metal2 ;
  RECT 673.440 46.820 674.560 50.060 ;
  LAYER metal1 ;
  RECT 673.440 46.820 674.560 50.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 38.980 674.560 42.220 ;
  LAYER metal4 ;
  RECT 673.440 38.980 674.560 42.220 ;
  LAYER metal3 ;
  RECT 673.440 38.980 674.560 42.220 ;
  LAYER metal2 ;
  RECT 673.440 38.980 674.560 42.220 ;
  LAYER metal1 ;
  RECT 673.440 38.980 674.560 42.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 31.140 674.560 34.380 ;
  LAYER metal4 ;
  RECT 673.440 31.140 674.560 34.380 ;
  LAYER metal3 ;
  RECT 673.440 31.140 674.560 34.380 ;
  LAYER metal2 ;
  RECT 673.440 31.140 674.560 34.380 ;
  LAYER metal1 ;
  RECT 673.440 31.140 674.560 34.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 23.300 674.560 26.540 ;
  LAYER metal4 ;
  RECT 673.440 23.300 674.560 26.540 ;
  LAYER metal3 ;
  RECT 673.440 23.300 674.560 26.540 ;
  LAYER metal2 ;
  RECT 673.440 23.300 674.560 26.540 ;
  LAYER metal1 ;
  RECT 673.440 23.300 674.560 26.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 15.460 674.560 18.700 ;
  LAYER metal4 ;
  RECT 673.440 15.460 674.560 18.700 ;
  LAYER metal3 ;
  RECT 673.440 15.460 674.560 18.700 ;
  LAYER metal2 ;
  RECT 673.440 15.460 674.560 18.700 ;
  LAYER metal1 ;
  RECT 673.440 15.460 674.560 18.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 7.620 674.560 10.860 ;
  LAYER metal4 ;
  RECT 673.440 7.620 674.560 10.860 ;
  LAYER metal3 ;
  RECT 673.440 7.620 674.560 10.860 ;
  LAYER metal2 ;
  RECT 673.440 7.620 674.560 10.860 ;
  LAYER metal1 ;
  RECT 673.440 7.620 674.560 10.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 634.820 1.120 638.060 ;
  LAYER metal4 ;
  RECT 0.000 634.820 1.120 638.060 ;
  LAYER metal3 ;
  RECT 0.000 634.820 1.120 638.060 ;
  LAYER metal2 ;
  RECT 0.000 634.820 1.120 638.060 ;
  LAYER metal1 ;
  RECT 0.000 634.820 1.120 638.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 595.620 1.120 598.860 ;
  LAYER metal4 ;
  RECT 0.000 595.620 1.120 598.860 ;
  LAYER metal3 ;
  RECT 0.000 595.620 1.120 598.860 ;
  LAYER metal2 ;
  RECT 0.000 595.620 1.120 598.860 ;
  LAYER metal1 ;
  RECT 0.000 595.620 1.120 598.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 587.780 1.120 591.020 ;
  LAYER metal4 ;
  RECT 0.000 587.780 1.120 591.020 ;
  LAYER metal3 ;
  RECT 0.000 587.780 1.120 591.020 ;
  LAYER metal2 ;
  RECT 0.000 587.780 1.120 591.020 ;
  LAYER metal1 ;
  RECT 0.000 587.780 1.120 591.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 579.940 1.120 583.180 ;
  LAYER metal4 ;
  RECT 0.000 579.940 1.120 583.180 ;
  LAYER metal3 ;
  RECT 0.000 579.940 1.120 583.180 ;
  LAYER metal2 ;
  RECT 0.000 579.940 1.120 583.180 ;
  LAYER metal1 ;
  RECT 0.000 579.940 1.120 583.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 572.100 1.120 575.340 ;
  LAYER metal4 ;
  RECT 0.000 572.100 1.120 575.340 ;
  LAYER metal3 ;
  RECT 0.000 572.100 1.120 575.340 ;
  LAYER metal2 ;
  RECT 0.000 572.100 1.120 575.340 ;
  LAYER metal1 ;
  RECT 0.000 572.100 1.120 575.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 564.260 1.120 567.500 ;
  LAYER metal4 ;
  RECT 0.000 564.260 1.120 567.500 ;
  LAYER metal3 ;
  RECT 0.000 564.260 1.120 567.500 ;
  LAYER metal2 ;
  RECT 0.000 564.260 1.120 567.500 ;
  LAYER metal1 ;
  RECT 0.000 564.260 1.120 567.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 556.420 1.120 559.660 ;
  LAYER metal4 ;
  RECT 0.000 556.420 1.120 559.660 ;
  LAYER metal3 ;
  RECT 0.000 556.420 1.120 559.660 ;
  LAYER metal2 ;
  RECT 0.000 556.420 1.120 559.660 ;
  LAYER metal1 ;
  RECT 0.000 556.420 1.120 559.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 517.220 1.120 520.460 ;
  LAYER metal4 ;
  RECT 0.000 517.220 1.120 520.460 ;
  LAYER metal3 ;
  RECT 0.000 517.220 1.120 520.460 ;
  LAYER metal2 ;
  RECT 0.000 517.220 1.120 520.460 ;
  LAYER metal1 ;
  RECT 0.000 517.220 1.120 520.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 509.380 1.120 512.620 ;
  LAYER metal4 ;
  RECT 0.000 509.380 1.120 512.620 ;
  LAYER metal3 ;
  RECT 0.000 509.380 1.120 512.620 ;
  LAYER metal2 ;
  RECT 0.000 509.380 1.120 512.620 ;
  LAYER metal1 ;
  RECT 0.000 509.380 1.120 512.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 501.540 1.120 504.780 ;
  LAYER metal4 ;
  RECT 0.000 501.540 1.120 504.780 ;
  LAYER metal3 ;
  RECT 0.000 501.540 1.120 504.780 ;
  LAYER metal2 ;
  RECT 0.000 501.540 1.120 504.780 ;
  LAYER metal1 ;
  RECT 0.000 501.540 1.120 504.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 493.700 1.120 496.940 ;
  LAYER metal4 ;
  RECT 0.000 493.700 1.120 496.940 ;
  LAYER metal3 ;
  RECT 0.000 493.700 1.120 496.940 ;
  LAYER metal2 ;
  RECT 0.000 493.700 1.120 496.940 ;
  LAYER metal1 ;
  RECT 0.000 493.700 1.120 496.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal4 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal3 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal2 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal1 ;
  RECT 0.000 485.860 1.120 489.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal4 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal3 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal2 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal1 ;
  RECT 0.000 478.020 1.120 481.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal4 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal3 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal2 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal1 ;
  RECT 0.000 438.820 1.120 442.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal4 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal3 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal2 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal1 ;
  RECT 0.000 430.980 1.120 434.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal4 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal3 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal2 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal1 ;
  RECT 0.000 423.140 1.120 426.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal4 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal3 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal2 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal1 ;
  RECT 0.000 415.300 1.120 418.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal4 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal3 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal2 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal1 ;
  RECT 0.000 407.460 1.120 410.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal4 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal3 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal2 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal1 ;
  RECT 0.000 399.620 1.120 402.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal4 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal3 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal2 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal1 ;
  RECT 0.000 360.420 1.120 363.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal4 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal3 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal2 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal1 ;
  RECT 0.000 352.580 1.120 355.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal4 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal3 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal2 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal1 ;
  RECT 0.000 344.740 1.120 347.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal4 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal3 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal2 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal1 ;
  RECT 0.000 336.900 1.120 340.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal4 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal3 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal2 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal1 ;
  RECT 0.000 329.060 1.120 332.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal4 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal3 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal2 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal1 ;
  RECT 0.000 321.220 1.120 324.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal4 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal3 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal2 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal1 ;
  RECT 0.000 282.020 1.120 285.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal4 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal3 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal2 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal1 ;
  RECT 0.000 274.180 1.120 277.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal4 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal3 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal2 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal1 ;
  RECT 0.000 266.340 1.120 269.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal4 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal3 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal2 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal1 ;
  RECT 0.000 258.500 1.120 261.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal4 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal3 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal2 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal1 ;
  RECT 0.000 250.660 1.120 253.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal4 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal3 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal2 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal1 ;
  RECT 0.000 242.820 1.120 246.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal4 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal3 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal2 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal1 ;
  RECT 0.000 203.620 1.120 206.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal4 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal3 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal2 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal1 ;
  RECT 0.000 195.780 1.120 199.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal4 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal3 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal2 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal1 ;
  RECT 0.000 187.940 1.120 191.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal4 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal3 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal2 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal1 ;
  RECT 0.000 180.100 1.120 183.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal4 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal3 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal2 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal1 ;
  RECT 0.000 172.260 1.120 175.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal4 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal3 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal2 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal1 ;
  RECT 0.000 164.420 1.120 167.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal4 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal3 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal2 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal1 ;
  RECT 0.000 125.220 1.120 128.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal4 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal3 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal2 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal1 ;
  RECT 0.000 117.380 1.120 120.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal4 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal3 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal2 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal1 ;
  RECT 0.000 109.540 1.120 112.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal4 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal3 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal2 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal1 ;
  RECT 0.000 101.700 1.120 104.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal4 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal3 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal2 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal1 ;
  RECT 0.000 93.860 1.120 97.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal4 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal3 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal2 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal1 ;
  RECT 0.000 86.020 1.120 89.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal4 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal3 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal2 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal1 ;
  RECT 0.000 46.820 1.120 50.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal4 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal3 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal2 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal1 ;
  RECT 0.000 38.980 1.120 42.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal4 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal3 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal2 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal1 ;
  RECT 0.000 31.140 1.120 34.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal4 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal3 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal2 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal1 ;
  RECT 0.000 23.300 1.120 26.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal4 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal3 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal2 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal1 ;
  RECT 0.000 15.460 1.120 18.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal4 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal3 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal2 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal1 ;
  RECT 0.000 7.620 1.120 10.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 644.580 646.800 648.120 647.920 ;
  LAYER metal4 ;
  RECT 644.580 646.800 648.120 647.920 ;
  LAYER metal3 ;
  RECT 644.580 646.800 648.120 647.920 ;
  LAYER metal2 ;
  RECT 644.580 646.800 648.120 647.920 ;
  LAYER metal1 ;
  RECT 644.580 646.800 648.120 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 631.560 646.800 635.100 647.920 ;
  LAYER metal4 ;
  RECT 631.560 646.800 635.100 647.920 ;
  LAYER metal3 ;
  RECT 631.560 646.800 635.100 647.920 ;
  LAYER metal2 ;
  RECT 631.560 646.800 635.100 647.920 ;
  LAYER metal1 ;
  RECT 631.560 646.800 635.100 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 617.920 646.800 621.460 647.920 ;
  LAYER metal4 ;
  RECT 617.920 646.800 621.460 647.920 ;
  LAYER metal3 ;
  RECT 617.920 646.800 621.460 647.920 ;
  LAYER metal2 ;
  RECT 617.920 646.800 621.460 647.920 ;
  LAYER metal1 ;
  RECT 617.920 646.800 621.460 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 604.280 646.800 607.820 647.920 ;
  LAYER metal4 ;
  RECT 604.280 646.800 607.820 647.920 ;
  LAYER metal3 ;
  RECT 604.280 646.800 607.820 647.920 ;
  LAYER metal2 ;
  RECT 604.280 646.800 607.820 647.920 ;
  LAYER metal1 ;
  RECT 604.280 646.800 607.820 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 591.260 646.800 594.800 647.920 ;
  LAYER metal4 ;
  RECT 591.260 646.800 594.800 647.920 ;
  LAYER metal3 ;
  RECT 591.260 646.800 594.800 647.920 ;
  LAYER metal2 ;
  RECT 591.260 646.800 594.800 647.920 ;
  LAYER metal1 ;
  RECT 591.260 646.800 594.800 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 577.620 646.800 581.160 647.920 ;
  LAYER metal4 ;
  RECT 577.620 646.800 581.160 647.920 ;
  LAYER metal3 ;
  RECT 577.620 646.800 581.160 647.920 ;
  LAYER metal2 ;
  RECT 577.620 646.800 581.160 647.920 ;
  LAYER metal1 ;
  RECT 577.620 646.800 581.160 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 510.660 646.800 514.200 647.920 ;
  LAYER metal4 ;
  RECT 510.660 646.800 514.200 647.920 ;
  LAYER metal3 ;
  RECT 510.660 646.800 514.200 647.920 ;
  LAYER metal2 ;
  RECT 510.660 646.800 514.200 647.920 ;
  LAYER metal1 ;
  RECT 510.660 646.800 514.200 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 497.020 646.800 500.560 647.920 ;
  LAYER metal4 ;
  RECT 497.020 646.800 500.560 647.920 ;
  LAYER metal3 ;
  RECT 497.020 646.800 500.560 647.920 ;
  LAYER metal2 ;
  RECT 497.020 646.800 500.560 647.920 ;
  LAYER metal1 ;
  RECT 497.020 646.800 500.560 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 483.380 646.800 486.920 647.920 ;
  LAYER metal4 ;
  RECT 483.380 646.800 486.920 647.920 ;
  LAYER metal3 ;
  RECT 483.380 646.800 486.920 647.920 ;
  LAYER metal2 ;
  RECT 483.380 646.800 486.920 647.920 ;
  LAYER metal1 ;
  RECT 483.380 646.800 486.920 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 469.740 646.800 473.280 647.920 ;
  LAYER metal4 ;
  RECT 469.740 646.800 473.280 647.920 ;
  LAYER metal3 ;
  RECT 469.740 646.800 473.280 647.920 ;
  LAYER metal2 ;
  RECT 469.740 646.800 473.280 647.920 ;
  LAYER metal1 ;
  RECT 469.740 646.800 473.280 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 456.720 646.800 460.260 647.920 ;
  LAYER metal4 ;
  RECT 456.720 646.800 460.260 647.920 ;
  LAYER metal3 ;
  RECT 456.720 646.800 460.260 647.920 ;
  LAYER metal2 ;
  RECT 456.720 646.800 460.260 647.920 ;
  LAYER metal1 ;
  RECT 456.720 646.800 460.260 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 443.080 646.800 446.620 647.920 ;
  LAYER metal4 ;
  RECT 443.080 646.800 446.620 647.920 ;
  LAYER metal3 ;
  RECT 443.080 646.800 446.620 647.920 ;
  LAYER metal2 ;
  RECT 443.080 646.800 446.620 647.920 ;
  LAYER metal1 ;
  RECT 443.080 646.800 446.620 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 381.080 646.800 384.620 647.920 ;
  LAYER metal4 ;
  RECT 381.080 646.800 384.620 647.920 ;
  LAYER metal3 ;
  RECT 381.080 646.800 384.620 647.920 ;
  LAYER metal2 ;
  RECT 381.080 646.800 384.620 647.920 ;
  LAYER metal1 ;
  RECT 381.080 646.800 384.620 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 352.560 646.800 356.100 647.920 ;
  LAYER metal4 ;
  RECT 352.560 646.800 356.100 647.920 ;
  LAYER metal3 ;
  RECT 352.560 646.800 356.100 647.920 ;
  LAYER metal2 ;
  RECT 352.560 646.800 356.100 647.920 ;
  LAYER metal1 ;
  RECT 352.560 646.800 356.100 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 328.380 646.800 331.920 647.920 ;
  LAYER metal4 ;
  RECT 328.380 646.800 331.920 647.920 ;
  LAYER metal3 ;
  RECT 328.380 646.800 331.920 647.920 ;
  LAYER metal2 ;
  RECT 328.380 646.800 331.920 647.920 ;
  LAYER metal1 ;
  RECT 328.380 646.800 331.920 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 302.340 646.800 305.880 647.920 ;
  LAYER metal4 ;
  RECT 302.340 646.800 305.880 647.920 ;
  LAYER metal3 ;
  RECT 302.340 646.800 305.880 647.920 ;
  LAYER metal2 ;
  RECT 302.340 646.800 305.880 647.920 ;
  LAYER metal1 ;
  RECT 302.340 646.800 305.880 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 283.120 646.800 286.660 647.920 ;
  LAYER metal4 ;
  RECT 283.120 646.800 286.660 647.920 ;
  LAYER metal3 ;
  RECT 283.120 646.800 286.660 647.920 ;
  LAYER metal2 ;
  RECT 283.120 646.800 286.660 647.920 ;
  LAYER metal1 ;
  RECT 283.120 646.800 286.660 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 274.440 646.800 277.980 647.920 ;
  LAYER metal4 ;
  RECT 274.440 646.800 277.980 647.920 ;
  LAYER metal3 ;
  RECT 274.440 646.800 277.980 647.920 ;
  LAYER metal2 ;
  RECT 274.440 646.800 277.980 647.920 ;
  LAYER metal1 ;
  RECT 274.440 646.800 277.980 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 207.480 646.800 211.020 647.920 ;
  LAYER metal4 ;
  RECT 207.480 646.800 211.020 647.920 ;
  LAYER metal3 ;
  RECT 207.480 646.800 211.020 647.920 ;
  LAYER metal2 ;
  RECT 207.480 646.800 211.020 647.920 ;
  LAYER metal1 ;
  RECT 207.480 646.800 211.020 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 193.840 646.800 197.380 647.920 ;
  LAYER metal4 ;
  RECT 193.840 646.800 197.380 647.920 ;
  LAYER metal3 ;
  RECT 193.840 646.800 197.380 647.920 ;
  LAYER metal2 ;
  RECT 193.840 646.800 197.380 647.920 ;
  LAYER metal1 ;
  RECT 193.840 646.800 197.380 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 180.820 646.800 184.360 647.920 ;
  LAYER metal4 ;
  RECT 180.820 646.800 184.360 647.920 ;
  LAYER metal3 ;
  RECT 180.820 646.800 184.360 647.920 ;
  LAYER metal2 ;
  RECT 180.820 646.800 184.360 647.920 ;
  LAYER metal1 ;
  RECT 180.820 646.800 184.360 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 167.180 646.800 170.720 647.920 ;
  LAYER metal4 ;
  RECT 167.180 646.800 170.720 647.920 ;
  LAYER metal3 ;
  RECT 167.180 646.800 170.720 647.920 ;
  LAYER metal2 ;
  RECT 167.180 646.800 170.720 647.920 ;
  LAYER metal1 ;
  RECT 167.180 646.800 170.720 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 153.540 646.800 157.080 647.920 ;
  LAYER metal4 ;
  RECT 153.540 646.800 157.080 647.920 ;
  LAYER metal3 ;
  RECT 153.540 646.800 157.080 647.920 ;
  LAYER metal2 ;
  RECT 153.540 646.800 157.080 647.920 ;
  LAYER metal1 ;
  RECT 153.540 646.800 157.080 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 140.520 646.800 144.060 647.920 ;
  LAYER metal4 ;
  RECT 140.520 646.800 144.060 647.920 ;
  LAYER metal3 ;
  RECT 140.520 646.800 144.060 647.920 ;
  LAYER metal2 ;
  RECT 140.520 646.800 144.060 647.920 ;
  LAYER metal1 ;
  RECT 140.520 646.800 144.060 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 72.940 646.800 76.480 647.920 ;
  LAYER metal4 ;
  RECT 72.940 646.800 76.480 647.920 ;
  LAYER metal3 ;
  RECT 72.940 646.800 76.480 647.920 ;
  LAYER metal2 ;
  RECT 72.940 646.800 76.480 647.920 ;
  LAYER metal1 ;
  RECT 72.940 646.800 76.480 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 59.300 646.800 62.840 647.920 ;
  LAYER metal4 ;
  RECT 59.300 646.800 62.840 647.920 ;
  LAYER metal3 ;
  RECT 59.300 646.800 62.840 647.920 ;
  LAYER metal2 ;
  RECT 59.300 646.800 62.840 647.920 ;
  LAYER metal1 ;
  RECT 59.300 646.800 62.840 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 46.280 646.800 49.820 647.920 ;
  LAYER metal4 ;
  RECT 46.280 646.800 49.820 647.920 ;
  LAYER metal3 ;
  RECT 46.280 646.800 49.820 647.920 ;
  LAYER metal2 ;
  RECT 46.280 646.800 49.820 647.920 ;
  LAYER metal1 ;
  RECT 46.280 646.800 49.820 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 32.640 646.800 36.180 647.920 ;
  LAYER metal4 ;
  RECT 32.640 646.800 36.180 647.920 ;
  LAYER metal3 ;
  RECT 32.640 646.800 36.180 647.920 ;
  LAYER metal2 ;
  RECT 32.640 646.800 36.180 647.920 ;
  LAYER metal1 ;
  RECT 32.640 646.800 36.180 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 19.000 646.800 22.540 647.920 ;
  LAYER metal4 ;
  RECT 19.000 646.800 22.540 647.920 ;
  LAYER metal3 ;
  RECT 19.000 646.800 22.540 647.920 ;
  LAYER metal2 ;
  RECT 19.000 646.800 22.540 647.920 ;
  LAYER metal1 ;
  RECT 19.000 646.800 22.540 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 7.220 646.800 10.760 647.920 ;
  LAYER metal4 ;
  RECT 7.220 646.800 10.760 647.920 ;
  LAYER metal3 ;
  RECT 7.220 646.800 10.760 647.920 ;
  LAYER metal2 ;
  RECT 7.220 646.800 10.760 647.920 ;
  LAYER metal1 ;
  RECT 7.220 646.800 10.760 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 644.580 0.000 648.120 1.120 ;
  LAYER metal4 ;
  RECT 644.580 0.000 648.120 1.120 ;
  LAYER metal3 ;
  RECT 644.580 0.000 648.120 1.120 ;
  LAYER metal2 ;
  RECT 644.580 0.000 648.120 1.120 ;
  LAYER metal1 ;
  RECT 644.580 0.000 648.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 631.560 0.000 635.100 1.120 ;
  LAYER metal4 ;
  RECT 631.560 0.000 635.100 1.120 ;
  LAYER metal3 ;
  RECT 631.560 0.000 635.100 1.120 ;
  LAYER metal2 ;
  RECT 631.560 0.000 635.100 1.120 ;
  LAYER metal1 ;
  RECT 631.560 0.000 635.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 617.920 0.000 621.460 1.120 ;
  LAYER metal4 ;
  RECT 617.920 0.000 621.460 1.120 ;
  LAYER metal3 ;
  RECT 617.920 0.000 621.460 1.120 ;
  LAYER metal2 ;
  RECT 617.920 0.000 621.460 1.120 ;
  LAYER metal1 ;
  RECT 617.920 0.000 621.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 604.280 0.000 607.820 1.120 ;
  LAYER metal4 ;
  RECT 604.280 0.000 607.820 1.120 ;
  LAYER metal3 ;
  RECT 604.280 0.000 607.820 1.120 ;
  LAYER metal2 ;
  RECT 604.280 0.000 607.820 1.120 ;
  LAYER metal1 ;
  RECT 604.280 0.000 607.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 591.260 0.000 594.800 1.120 ;
  LAYER metal4 ;
  RECT 591.260 0.000 594.800 1.120 ;
  LAYER metal3 ;
  RECT 591.260 0.000 594.800 1.120 ;
  LAYER metal2 ;
  RECT 591.260 0.000 594.800 1.120 ;
  LAYER metal1 ;
  RECT 591.260 0.000 594.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 577.620 0.000 581.160 1.120 ;
  LAYER metal4 ;
  RECT 577.620 0.000 581.160 1.120 ;
  LAYER metal3 ;
  RECT 577.620 0.000 581.160 1.120 ;
  LAYER metal2 ;
  RECT 577.620 0.000 581.160 1.120 ;
  LAYER metal1 ;
  RECT 577.620 0.000 581.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 510.660 0.000 514.200 1.120 ;
  LAYER metal4 ;
  RECT 510.660 0.000 514.200 1.120 ;
  LAYER metal3 ;
  RECT 510.660 0.000 514.200 1.120 ;
  LAYER metal2 ;
  RECT 510.660 0.000 514.200 1.120 ;
  LAYER metal1 ;
  RECT 510.660 0.000 514.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 497.020 0.000 500.560 1.120 ;
  LAYER metal4 ;
  RECT 497.020 0.000 500.560 1.120 ;
  LAYER metal3 ;
  RECT 497.020 0.000 500.560 1.120 ;
  LAYER metal2 ;
  RECT 497.020 0.000 500.560 1.120 ;
  LAYER metal1 ;
  RECT 497.020 0.000 500.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 483.380 0.000 486.920 1.120 ;
  LAYER metal4 ;
  RECT 483.380 0.000 486.920 1.120 ;
  LAYER metal3 ;
  RECT 483.380 0.000 486.920 1.120 ;
  LAYER metal2 ;
  RECT 483.380 0.000 486.920 1.120 ;
  LAYER metal1 ;
  RECT 483.380 0.000 486.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 469.740 0.000 473.280 1.120 ;
  LAYER metal4 ;
  RECT 469.740 0.000 473.280 1.120 ;
  LAYER metal3 ;
  RECT 469.740 0.000 473.280 1.120 ;
  LAYER metal2 ;
  RECT 469.740 0.000 473.280 1.120 ;
  LAYER metal1 ;
  RECT 469.740 0.000 473.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 456.720 0.000 460.260 1.120 ;
  LAYER metal4 ;
  RECT 456.720 0.000 460.260 1.120 ;
  LAYER metal3 ;
  RECT 456.720 0.000 460.260 1.120 ;
  LAYER metal2 ;
  RECT 456.720 0.000 460.260 1.120 ;
  LAYER metal1 ;
  RECT 456.720 0.000 460.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 443.080 0.000 446.620 1.120 ;
  LAYER metal4 ;
  RECT 443.080 0.000 446.620 1.120 ;
  LAYER metal3 ;
  RECT 443.080 0.000 446.620 1.120 ;
  LAYER metal2 ;
  RECT 443.080 0.000 446.620 1.120 ;
  LAYER metal1 ;
  RECT 443.080 0.000 446.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 381.080 0.000 384.620 1.120 ;
  LAYER metal4 ;
  RECT 381.080 0.000 384.620 1.120 ;
  LAYER metal3 ;
  RECT 381.080 0.000 384.620 1.120 ;
  LAYER metal2 ;
  RECT 381.080 0.000 384.620 1.120 ;
  LAYER metal1 ;
  RECT 381.080 0.000 384.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 352.560 0.000 356.100 1.120 ;
  LAYER metal4 ;
  RECT 352.560 0.000 356.100 1.120 ;
  LAYER metal3 ;
  RECT 352.560 0.000 356.100 1.120 ;
  LAYER metal2 ;
  RECT 352.560 0.000 356.100 1.120 ;
  LAYER metal1 ;
  RECT 352.560 0.000 356.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal4 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal3 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal2 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal1 ;
  RECT 328.380 0.000 331.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 302.340 0.000 305.880 1.120 ;
  LAYER metal4 ;
  RECT 302.340 0.000 305.880 1.120 ;
  LAYER metal3 ;
  RECT 302.340 0.000 305.880 1.120 ;
  LAYER metal2 ;
  RECT 302.340 0.000 305.880 1.120 ;
  LAYER metal1 ;
  RECT 302.340 0.000 305.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal4 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal3 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal2 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal1 ;
  RECT 283.120 0.000 286.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal4 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal3 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal2 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal1 ;
  RECT 274.440 0.000 277.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal4 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal3 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal2 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal1 ;
  RECT 207.480 0.000 211.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal4 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal3 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal2 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal1 ;
  RECT 193.840 0.000 197.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal4 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal3 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal2 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal1 ;
  RECT 180.820 0.000 184.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal4 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal3 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal2 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal1 ;
  RECT 167.180 0.000 170.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal4 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal3 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal2 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal1 ;
  RECT 153.540 0.000 157.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal4 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal3 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal2 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal1 ;
  RECT 140.520 0.000 144.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal4 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal3 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal2 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal1 ;
  RECT 72.940 0.000 76.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal4 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal3 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal2 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal1 ;
  RECT 59.300 0.000 62.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal4 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal3 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal2 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal1 ;
  RECT 46.280 0.000 49.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal4 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal3 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal2 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal1 ;
  RECT 32.640 0.000 36.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal4 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal3 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal2 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal1 ;
  RECT 19.000 0.000 22.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal4 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal3 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal2 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal1 ;
  RECT 7.220 0.000 10.760 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal5 ;
  RECT 673.440 599.540 674.560 602.780 ;
  LAYER metal4 ;
  RECT 673.440 599.540 674.560 602.780 ;
  LAYER metal3 ;
  RECT 673.440 599.540 674.560 602.780 ;
  LAYER metal2 ;
  RECT 673.440 599.540 674.560 602.780 ;
  LAYER metal1 ;
  RECT 673.440 599.540 674.560 602.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 591.700 674.560 594.940 ;
  LAYER metal4 ;
  RECT 673.440 591.700 674.560 594.940 ;
  LAYER metal3 ;
  RECT 673.440 591.700 674.560 594.940 ;
  LAYER metal2 ;
  RECT 673.440 591.700 674.560 594.940 ;
  LAYER metal1 ;
  RECT 673.440 591.700 674.560 594.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 583.860 674.560 587.100 ;
  LAYER metal4 ;
  RECT 673.440 583.860 674.560 587.100 ;
  LAYER metal3 ;
  RECT 673.440 583.860 674.560 587.100 ;
  LAYER metal2 ;
  RECT 673.440 583.860 674.560 587.100 ;
  LAYER metal1 ;
  RECT 673.440 583.860 674.560 587.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 576.020 674.560 579.260 ;
  LAYER metal4 ;
  RECT 673.440 576.020 674.560 579.260 ;
  LAYER metal3 ;
  RECT 673.440 576.020 674.560 579.260 ;
  LAYER metal2 ;
  RECT 673.440 576.020 674.560 579.260 ;
  LAYER metal1 ;
  RECT 673.440 576.020 674.560 579.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 568.180 674.560 571.420 ;
  LAYER metal4 ;
  RECT 673.440 568.180 674.560 571.420 ;
  LAYER metal3 ;
  RECT 673.440 568.180 674.560 571.420 ;
  LAYER metal2 ;
  RECT 673.440 568.180 674.560 571.420 ;
  LAYER metal1 ;
  RECT 673.440 568.180 674.560 571.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 560.340 674.560 563.580 ;
  LAYER metal4 ;
  RECT 673.440 560.340 674.560 563.580 ;
  LAYER metal3 ;
  RECT 673.440 560.340 674.560 563.580 ;
  LAYER metal2 ;
  RECT 673.440 560.340 674.560 563.580 ;
  LAYER metal1 ;
  RECT 673.440 560.340 674.560 563.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 521.140 674.560 524.380 ;
  LAYER metal4 ;
  RECT 673.440 521.140 674.560 524.380 ;
  LAYER metal3 ;
  RECT 673.440 521.140 674.560 524.380 ;
  LAYER metal2 ;
  RECT 673.440 521.140 674.560 524.380 ;
  LAYER metal1 ;
  RECT 673.440 521.140 674.560 524.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 513.300 674.560 516.540 ;
  LAYER metal4 ;
  RECT 673.440 513.300 674.560 516.540 ;
  LAYER metal3 ;
  RECT 673.440 513.300 674.560 516.540 ;
  LAYER metal2 ;
  RECT 673.440 513.300 674.560 516.540 ;
  LAYER metal1 ;
  RECT 673.440 513.300 674.560 516.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 505.460 674.560 508.700 ;
  LAYER metal4 ;
  RECT 673.440 505.460 674.560 508.700 ;
  LAYER metal3 ;
  RECT 673.440 505.460 674.560 508.700 ;
  LAYER metal2 ;
  RECT 673.440 505.460 674.560 508.700 ;
  LAYER metal1 ;
  RECT 673.440 505.460 674.560 508.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 497.620 674.560 500.860 ;
  LAYER metal4 ;
  RECT 673.440 497.620 674.560 500.860 ;
  LAYER metal3 ;
  RECT 673.440 497.620 674.560 500.860 ;
  LAYER metal2 ;
  RECT 673.440 497.620 674.560 500.860 ;
  LAYER metal1 ;
  RECT 673.440 497.620 674.560 500.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 489.780 674.560 493.020 ;
  LAYER metal4 ;
  RECT 673.440 489.780 674.560 493.020 ;
  LAYER metal3 ;
  RECT 673.440 489.780 674.560 493.020 ;
  LAYER metal2 ;
  RECT 673.440 489.780 674.560 493.020 ;
  LAYER metal1 ;
  RECT 673.440 489.780 674.560 493.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 481.940 674.560 485.180 ;
  LAYER metal4 ;
  RECT 673.440 481.940 674.560 485.180 ;
  LAYER metal3 ;
  RECT 673.440 481.940 674.560 485.180 ;
  LAYER metal2 ;
  RECT 673.440 481.940 674.560 485.180 ;
  LAYER metal1 ;
  RECT 673.440 481.940 674.560 485.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 442.740 674.560 445.980 ;
  LAYER metal4 ;
  RECT 673.440 442.740 674.560 445.980 ;
  LAYER metal3 ;
  RECT 673.440 442.740 674.560 445.980 ;
  LAYER metal2 ;
  RECT 673.440 442.740 674.560 445.980 ;
  LAYER metal1 ;
  RECT 673.440 442.740 674.560 445.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 434.900 674.560 438.140 ;
  LAYER metal4 ;
  RECT 673.440 434.900 674.560 438.140 ;
  LAYER metal3 ;
  RECT 673.440 434.900 674.560 438.140 ;
  LAYER metal2 ;
  RECT 673.440 434.900 674.560 438.140 ;
  LAYER metal1 ;
  RECT 673.440 434.900 674.560 438.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 427.060 674.560 430.300 ;
  LAYER metal4 ;
  RECT 673.440 427.060 674.560 430.300 ;
  LAYER metal3 ;
  RECT 673.440 427.060 674.560 430.300 ;
  LAYER metal2 ;
  RECT 673.440 427.060 674.560 430.300 ;
  LAYER metal1 ;
  RECT 673.440 427.060 674.560 430.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 419.220 674.560 422.460 ;
  LAYER metal4 ;
  RECT 673.440 419.220 674.560 422.460 ;
  LAYER metal3 ;
  RECT 673.440 419.220 674.560 422.460 ;
  LAYER metal2 ;
  RECT 673.440 419.220 674.560 422.460 ;
  LAYER metal1 ;
  RECT 673.440 419.220 674.560 422.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 411.380 674.560 414.620 ;
  LAYER metal4 ;
  RECT 673.440 411.380 674.560 414.620 ;
  LAYER metal3 ;
  RECT 673.440 411.380 674.560 414.620 ;
  LAYER metal2 ;
  RECT 673.440 411.380 674.560 414.620 ;
  LAYER metal1 ;
  RECT 673.440 411.380 674.560 414.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 403.540 674.560 406.780 ;
  LAYER metal4 ;
  RECT 673.440 403.540 674.560 406.780 ;
  LAYER metal3 ;
  RECT 673.440 403.540 674.560 406.780 ;
  LAYER metal2 ;
  RECT 673.440 403.540 674.560 406.780 ;
  LAYER metal1 ;
  RECT 673.440 403.540 674.560 406.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 364.340 674.560 367.580 ;
  LAYER metal4 ;
  RECT 673.440 364.340 674.560 367.580 ;
  LAYER metal3 ;
  RECT 673.440 364.340 674.560 367.580 ;
  LAYER metal2 ;
  RECT 673.440 364.340 674.560 367.580 ;
  LAYER metal1 ;
  RECT 673.440 364.340 674.560 367.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 356.500 674.560 359.740 ;
  LAYER metal4 ;
  RECT 673.440 356.500 674.560 359.740 ;
  LAYER metal3 ;
  RECT 673.440 356.500 674.560 359.740 ;
  LAYER metal2 ;
  RECT 673.440 356.500 674.560 359.740 ;
  LAYER metal1 ;
  RECT 673.440 356.500 674.560 359.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 348.660 674.560 351.900 ;
  LAYER metal4 ;
  RECT 673.440 348.660 674.560 351.900 ;
  LAYER metal3 ;
  RECT 673.440 348.660 674.560 351.900 ;
  LAYER metal2 ;
  RECT 673.440 348.660 674.560 351.900 ;
  LAYER metal1 ;
  RECT 673.440 348.660 674.560 351.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 340.820 674.560 344.060 ;
  LAYER metal4 ;
  RECT 673.440 340.820 674.560 344.060 ;
  LAYER metal3 ;
  RECT 673.440 340.820 674.560 344.060 ;
  LAYER metal2 ;
  RECT 673.440 340.820 674.560 344.060 ;
  LAYER metal1 ;
  RECT 673.440 340.820 674.560 344.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 332.980 674.560 336.220 ;
  LAYER metal4 ;
  RECT 673.440 332.980 674.560 336.220 ;
  LAYER metal3 ;
  RECT 673.440 332.980 674.560 336.220 ;
  LAYER metal2 ;
  RECT 673.440 332.980 674.560 336.220 ;
  LAYER metal1 ;
  RECT 673.440 332.980 674.560 336.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 325.140 674.560 328.380 ;
  LAYER metal4 ;
  RECT 673.440 325.140 674.560 328.380 ;
  LAYER metal3 ;
  RECT 673.440 325.140 674.560 328.380 ;
  LAYER metal2 ;
  RECT 673.440 325.140 674.560 328.380 ;
  LAYER metal1 ;
  RECT 673.440 325.140 674.560 328.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 285.940 674.560 289.180 ;
  LAYER metal4 ;
  RECT 673.440 285.940 674.560 289.180 ;
  LAYER metal3 ;
  RECT 673.440 285.940 674.560 289.180 ;
  LAYER metal2 ;
  RECT 673.440 285.940 674.560 289.180 ;
  LAYER metal1 ;
  RECT 673.440 285.940 674.560 289.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 278.100 674.560 281.340 ;
  LAYER metal4 ;
  RECT 673.440 278.100 674.560 281.340 ;
  LAYER metal3 ;
  RECT 673.440 278.100 674.560 281.340 ;
  LAYER metal2 ;
  RECT 673.440 278.100 674.560 281.340 ;
  LAYER metal1 ;
  RECT 673.440 278.100 674.560 281.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 270.260 674.560 273.500 ;
  LAYER metal4 ;
  RECT 673.440 270.260 674.560 273.500 ;
  LAYER metal3 ;
  RECT 673.440 270.260 674.560 273.500 ;
  LAYER metal2 ;
  RECT 673.440 270.260 674.560 273.500 ;
  LAYER metal1 ;
  RECT 673.440 270.260 674.560 273.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 262.420 674.560 265.660 ;
  LAYER metal4 ;
  RECT 673.440 262.420 674.560 265.660 ;
  LAYER metal3 ;
  RECT 673.440 262.420 674.560 265.660 ;
  LAYER metal2 ;
  RECT 673.440 262.420 674.560 265.660 ;
  LAYER metal1 ;
  RECT 673.440 262.420 674.560 265.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 254.580 674.560 257.820 ;
  LAYER metal4 ;
  RECT 673.440 254.580 674.560 257.820 ;
  LAYER metal3 ;
  RECT 673.440 254.580 674.560 257.820 ;
  LAYER metal2 ;
  RECT 673.440 254.580 674.560 257.820 ;
  LAYER metal1 ;
  RECT 673.440 254.580 674.560 257.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 246.740 674.560 249.980 ;
  LAYER metal4 ;
  RECT 673.440 246.740 674.560 249.980 ;
  LAYER metal3 ;
  RECT 673.440 246.740 674.560 249.980 ;
  LAYER metal2 ;
  RECT 673.440 246.740 674.560 249.980 ;
  LAYER metal1 ;
  RECT 673.440 246.740 674.560 249.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 207.540 674.560 210.780 ;
  LAYER metal4 ;
  RECT 673.440 207.540 674.560 210.780 ;
  LAYER metal3 ;
  RECT 673.440 207.540 674.560 210.780 ;
  LAYER metal2 ;
  RECT 673.440 207.540 674.560 210.780 ;
  LAYER metal1 ;
  RECT 673.440 207.540 674.560 210.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 199.700 674.560 202.940 ;
  LAYER metal4 ;
  RECT 673.440 199.700 674.560 202.940 ;
  LAYER metal3 ;
  RECT 673.440 199.700 674.560 202.940 ;
  LAYER metal2 ;
  RECT 673.440 199.700 674.560 202.940 ;
  LAYER metal1 ;
  RECT 673.440 199.700 674.560 202.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 191.860 674.560 195.100 ;
  LAYER metal4 ;
  RECT 673.440 191.860 674.560 195.100 ;
  LAYER metal3 ;
  RECT 673.440 191.860 674.560 195.100 ;
  LAYER metal2 ;
  RECT 673.440 191.860 674.560 195.100 ;
  LAYER metal1 ;
  RECT 673.440 191.860 674.560 195.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 184.020 674.560 187.260 ;
  LAYER metal4 ;
  RECT 673.440 184.020 674.560 187.260 ;
  LAYER metal3 ;
  RECT 673.440 184.020 674.560 187.260 ;
  LAYER metal2 ;
  RECT 673.440 184.020 674.560 187.260 ;
  LAYER metal1 ;
  RECT 673.440 184.020 674.560 187.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 176.180 674.560 179.420 ;
  LAYER metal4 ;
  RECT 673.440 176.180 674.560 179.420 ;
  LAYER metal3 ;
  RECT 673.440 176.180 674.560 179.420 ;
  LAYER metal2 ;
  RECT 673.440 176.180 674.560 179.420 ;
  LAYER metal1 ;
  RECT 673.440 176.180 674.560 179.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 168.340 674.560 171.580 ;
  LAYER metal4 ;
  RECT 673.440 168.340 674.560 171.580 ;
  LAYER metal3 ;
  RECT 673.440 168.340 674.560 171.580 ;
  LAYER metal2 ;
  RECT 673.440 168.340 674.560 171.580 ;
  LAYER metal1 ;
  RECT 673.440 168.340 674.560 171.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 129.140 674.560 132.380 ;
  LAYER metal4 ;
  RECT 673.440 129.140 674.560 132.380 ;
  LAYER metal3 ;
  RECT 673.440 129.140 674.560 132.380 ;
  LAYER metal2 ;
  RECT 673.440 129.140 674.560 132.380 ;
  LAYER metal1 ;
  RECT 673.440 129.140 674.560 132.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 121.300 674.560 124.540 ;
  LAYER metal4 ;
  RECT 673.440 121.300 674.560 124.540 ;
  LAYER metal3 ;
  RECT 673.440 121.300 674.560 124.540 ;
  LAYER metal2 ;
  RECT 673.440 121.300 674.560 124.540 ;
  LAYER metal1 ;
  RECT 673.440 121.300 674.560 124.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 113.460 674.560 116.700 ;
  LAYER metal4 ;
  RECT 673.440 113.460 674.560 116.700 ;
  LAYER metal3 ;
  RECT 673.440 113.460 674.560 116.700 ;
  LAYER metal2 ;
  RECT 673.440 113.460 674.560 116.700 ;
  LAYER metal1 ;
  RECT 673.440 113.460 674.560 116.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 105.620 674.560 108.860 ;
  LAYER metal4 ;
  RECT 673.440 105.620 674.560 108.860 ;
  LAYER metal3 ;
  RECT 673.440 105.620 674.560 108.860 ;
  LAYER metal2 ;
  RECT 673.440 105.620 674.560 108.860 ;
  LAYER metal1 ;
  RECT 673.440 105.620 674.560 108.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 97.780 674.560 101.020 ;
  LAYER metal4 ;
  RECT 673.440 97.780 674.560 101.020 ;
  LAYER metal3 ;
  RECT 673.440 97.780 674.560 101.020 ;
  LAYER metal2 ;
  RECT 673.440 97.780 674.560 101.020 ;
  LAYER metal1 ;
  RECT 673.440 97.780 674.560 101.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 89.940 674.560 93.180 ;
  LAYER metal4 ;
  RECT 673.440 89.940 674.560 93.180 ;
  LAYER metal3 ;
  RECT 673.440 89.940 674.560 93.180 ;
  LAYER metal2 ;
  RECT 673.440 89.940 674.560 93.180 ;
  LAYER metal1 ;
  RECT 673.440 89.940 674.560 93.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 50.740 674.560 53.980 ;
  LAYER metal4 ;
  RECT 673.440 50.740 674.560 53.980 ;
  LAYER metal3 ;
  RECT 673.440 50.740 674.560 53.980 ;
  LAYER metal2 ;
  RECT 673.440 50.740 674.560 53.980 ;
  LAYER metal1 ;
  RECT 673.440 50.740 674.560 53.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 42.900 674.560 46.140 ;
  LAYER metal4 ;
  RECT 673.440 42.900 674.560 46.140 ;
  LAYER metal3 ;
  RECT 673.440 42.900 674.560 46.140 ;
  LAYER metal2 ;
  RECT 673.440 42.900 674.560 46.140 ;
  LAYER metal1 ;
  RECT 673.440 42.900 674.560 46.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 35.060 674.560 38.300 ;
  LAYER metal4 ;
  RECT 673.440 35.060 674.560 38.300 ;
  LAYER metal3 ;
  RECT 673.440 35.060 674.560 38.300 ;
  LAYER metal2 ;
  RECT 673.440 35.060 674.560 38.300 ;
  LAYER metal1 ;
  RECT 673.440 35.060 674.560 38.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 27.220 674.560 30.460 ;
  LAYER metal4 ;
  RECT 673.440 27.220 674.560 30.460 ;
  LAYER metal3 ;
  RECT 673.440 27.220 674.560 30.460 ;
  LAYER metal2 ;
  RECT 673.440 27.220 674.560 30.460 ;
  LAYER metal1 ;
  RECT 673.440 27.220 674.560 30.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 19.380 674.560 22.620 ;
  LAYER metal4 ;
  RECT 673.440 19.380 674.560 22.620 ;
  LAYER metal3 ;
  RECT 673.440 19.380 674.560 22.620 ;
  LAYER metal2 ;
  RECT 673.440 19.380 674.560 22.620 ;
  LAYER metal1 ;
  RECT 673.440 19.380 674.560 22.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 673.440 11.540 674.560 14.780 ;
  LAYER metal4 ;
  RECT 673.440 11.540 674.560 14.780 ;
  LAYER metal3 ;
  RECT 673.440 11.540 674.560 14.780 ;
  LAYER metal2 ;
  RECT 673.440 11.540 674.560 14.780 ;
  LAYER metal1 ;
  RECT 673.440 11.540 674.560 14.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 599.540 1.120 602.780 ;
  LAYER metal4 ;
  RECT 0.000 599.540 1.120 602.780 ;
  LAYER metal3 ;
  RECT 0.000 599.540 1.120 602.780 ;
  LAYER metal2 ;
  RECT 0.000 599.540 1.120 602.780 ;
  LAYER metal1 ;
  RECT 0.000 599.540 1.120 602.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 591.700 1.120 594.940 ;
  LAYER metal4 ;
  RECT 0.000 591.700 1.120 594.940 ;
  LAYER metal3 ;
  RECT 0.000 591.700 1.120 594.940 ;
  LAYER metal2 ;
  RECT 0.000 591.700 1.120 594.940 ;
  LAYER metal1 ;
  RECT 0.000 591.700 1.120 594.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 583.860 1.120 587.100 ;
  LAYER metal4 ;
  RECT 0.000 583.860 1.120 587.100 ;
  LAYER metal3 ;
  RECT 0.000 583.860 1.120 587.100 ;
  LAYER metal2 ;
  RECT 0.000 583.860 1.120 587.100 ;
  LAYER metal1 ;
  RECT 0.000 583.860 1.120 587.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 576.020 1.120 579.260 ;
  LAYER metal4 ;
  RECT 0.000 576.020 1.120 579.260 ;
  LAYER metal3 ;
  RECT 0.000 576.020 1.120 579.260 ;
  LAYER metal2 ;
  RECT 0.000 576.020 1.120 579.260 ;
  LAYER metal1 ;
  RECT 0.000 576.020 1.120 579.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 568.180 1.120 571.420 ;
  LAYER metal4 ;
  RECT 0.000 568.180 1.120 571.420 ;
  LAYER metal3 ;
  RECT 0.000 568.180 1.120 571.420 ;
  LAYER metal2 ;
  RECT 0.000 568.180 1.120 571.420 ;
  LAYER metal1 ;
  RECT 0.000 568.180 1.120 571.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 560.340 1.120 563.580 ;
  LAYER metal4 ;
  RECT 0.000 560.340 1.120 563.580 ;
  LAYER metal3 ;
  RECT 0.000 560.340 1.120 563.580 ;
  LAYER metal2 ;
  RECT 0.000 560.340 1.120 563.580 ;
  LAYER metal1 ;
  RECT 0.000 560.340 1.120 563.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 521.140 1.120 524.380 ;
  LAYER metal4 ;
  RECT 0.000 521.140 1.120 524.380 ;
  LAYER metal3 ;
  RECT 0.000 521.140 1.120 524.380 ;
  LAYER metal2 ;
  RECT 0.000 521.140 1.120 524.380 ;
  LAYER metal1 ;
  RECT 0.000 521.140 1.120 524.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 513.300 1.120 516.540 ;
  LAYER metal4 ;
  RECT 0.000 513.300 1.120 516.540 ;
  LAYER metal3 ;
  RECT 0.000 513.300 1.120 516.540 ;
  LAYER metal2 ;
  RECT 0.000 513.300 1.120 516.540 ;
  LAYER metal1 ;
  RECT 0.000 513.300 1.120 516.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 505.460 1.120 508.700 ;
  LAYER metal4 ;
  RECT 0.000 505.460 1.120 508.700 ;
  LAYER metal3 ;
  RECT 0.000 505.460 1.120 508.700 ;
  LAYER metal2 ;
  RECT 0.000 505.460 1.120 508.700 ;
  LAYER metal1 ;
  RECT 0.000 505.460 1.120 508.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 497.620 1.120 500.860 ;
  LAYER metal4 ;
  RECT 0.000 497.620 1.120 500.860 ;
  LAYER metal3 ;
  RECT 0.000 497.620 1.120 500.860 ;
  LAYER metal2 ;
  RECT 0.000 497.620 1.120 500.860 ;
  LAYER metal1 ;
  RECT 0.000 497.620 1.120 500.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal4 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal3 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal2 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal1 ;
  RECT 0.000 489.780 1.120 493.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal4 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal3 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal2 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal1 ;
  RECT 0.000 481.940 1.120 485.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal4 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal3 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal2 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal1 ;
  RECT 0.000 442.740 1.120 445.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal4 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal3 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal2 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal1 ;
  RECT 0.000 434.900 1.120 438.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal4 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal3 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal2 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal1 ;
  RECT 0.000 427.060 1.120 430.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal4 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal3 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal2 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal1 ;
  RECT 0.000 419.220 1.120 422.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal4 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal3 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal2 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal1 ;
  RECT 0.000 411.380 1.120 414.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal4 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal3 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal2 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal1 ;
  RECT 0.000 403.540 1.120 406.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal4 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal3 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal2 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal1 ;
  RECT 0.000 364.340 1.120 367.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal4 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal3 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal2 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal1 ;
  RECT 0.000 356.500 1.120 359.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal4 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal3 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal2 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal1 ;
  RECT 0.000 348.660 1.120 351.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal4 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal3 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal2 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal1 ;
  RECT 0.000 340.820 1.120 344.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal4 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal3 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal2 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal1 ;
  RECT 0.000 332.980 1.120 336.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal4 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal3 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal2 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal1 ;
  RECT 0.000 325.140 1.120 328.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal4 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal3 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal2 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal1 ;
  RECT 0.000 285.940 1.120 289.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal4 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal3 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal2 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal1 ;
  RECT 0.000 278.100 1.120 281.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal4 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal3 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal2 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal1 ;
  RECT 0.000 270.260 1.120 273.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal4 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal3 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal2 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal1 ;
  RECT 0.000 262.420 1.120 265.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal4 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal3 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal2 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal1 ;
  RECT 0.000 254.580 1.120 257.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal4 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal3 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal2 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal1 ;
  RECT 0.000 246.740 1.120 249.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal4 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal3 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal2 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal1 ;
  RECT 0.000 207.540 1.120 210.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal4 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal3 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal2 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal1 ;
  RECT 0.000 199.700 1.120 202.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal4 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal3 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal2 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal1 ;
  RECT 0.000 191.860 1.120 195.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal4 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal3 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal2 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal1 ;
  RECT 0.000 184.020 1.120 187.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal4 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal3 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal2 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal1 ;
  RECT 0.000 176.180 1.120 179.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal4 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal3 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal2 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal1 ;
  RECT 0.000 168.340 1.120 171.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal4 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal3 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal2 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal1 ;
  RECT 0.000 129.140 1.120 132.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal4 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal3 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal2 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal1 ;
  RECT 0.000 121.300 1.120 124.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal4 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal3 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal2 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal1 ;
  RECT 0.000 113.460 1.120 116.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal4 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal3 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal2 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal1 ;
  RECT 0.000 105.620 1.120 108.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal4 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal3 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal2 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal1 ;
  RECT 0.000 97.780 1.120 101.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal4 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal3 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal2 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal1 ;
  RECT 0.000 89.940 1.120 93.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal4 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal3 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal2 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal1 ;
  RECT 0.000 50.740 1.120 53.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal4 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal3 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal2 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal1 ;
  RECT 0.000 42.900 1.120 46.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal4 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal3 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal2 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal1 ;
  RECT 0.000 35.060 1.120 38.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal4 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal3 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal2 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal1 ;
  RECT 0.000 27.220 1.120 30.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal4 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal3 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal2 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal1 ;
  RECT 0.000 19.380 1.120 22.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal4 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal3 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal2 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal1 ;
  RECT 0.000 11.540 1.120 14.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 653.880 646.800 657.420 647.920 ;
  LAYER metal4 ;
  RECT 653.880 646.800 657.420 647.920 ;
  LAYER metal3 ;
  RECT 653.880 646.800 657.420 647.920 ;
  LAYER metal2 ;
  RECT 653.880 646.800 657.420 647.920 ;
  LAYER metal1 ;
  RECT 653.880 646.800 657.420 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 640.240 646.800 643.780 647.920 ;
  LAYER metal4 ;
  RECT 640.240 646.800 643.780 647.920 ;
  LAYER metal3 ;
  RECT 640.240 646.800 643.780 647.920 ;
  LAYER metal2 ;
  RECT 640.240 646.800 643.780 647.920 ;
  LAYER metal1 ;
  RECT 640.240 646.800 643.780 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 627.220 646.800 630.760 647.920 ;
  LAYER metal4 ;
  RECT 627.220 646.800 630.760 647.920 ;
  LAYER metal3 ;
  RECT 627.220 646.800 630.760 647.920 ;
  LAYER metal2 ;
  RECT 627.220 646.800 630.760 647.920 ;
  LAYER metal1 ;
  RECT 627.220 646.800 630.760 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 613.580 646.800 617.120 647.920 ;
  LAYER metal4 ;
  RECT 613.580 646.800 617.120 647.920 ;
  LAYER metal3 ;
  RECT 613.580 646.800 617.120 647.920 ;
  LAYER metal2 ;
  RECT 613.580 646.800 617.120 647.920 ;
  LAYER metal1 ;
  RECT 613.580 646.800 617.120 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 599.940 646.800 603.480 647.920 ;
  LAYER metal4 ;
  RECT 599.940 646.800 603.480 647.920 ;
  LAYER metal3 ;
  RECT 599.940 646.800 603.480 647.920 ;
  LAYER metal2 ;
  RECT 599.940 646.800 603.480 647.920 ;
  LAYER metal1 ;
  RECT 599.940 646.800 603.480 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 586.920 646.800 590.460 647.920 ;
  LAYER metal4 ;
  RECT 586.920 646.800 590.460 647.920 ;
  LAYER metal3 ;
  RECT 586.920 646.800 590.460 647.920 ;
  LAYER metal2 ;
  RECT 586.920 646.800 590.460 647.920 ;
  LAYER metal1 ;
  RECT 586.920 646.800 590.460 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 519.340 646.800 522.880 647.920 ;
  LAYER metal4 ;
  RECT 519.340 646.800 522.880 647.920 ;
  LAYER metal3 ;
  RECT 519.340 646.800 522.880 647.920 ;
  LAYER metal2 ;
  RECT 519.340 646.800 522.880 647.920 ;
  LAYER metal1 ;
  RECT 519.340 646.800 522.880 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 506.320 646.800 509.860 647.920 ;
  LAYER metal4 ;
  RECT 506.320 646.800 509.860 647.920 ;
  LAYER metal3 ;
  RECT 506.320 646.800 509.860 647.920 ;
  LAYER metal2 ;
  RECT 506.320 646.800 509.860 647.920 ;
  LAYER metal1 ;
  RECT 506.320 646.800 509.860 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 492.680 646.800 496.220 647.920 ;
  LAYER metal4 ;
  RECT 492.680 646.800 496.220 647.920 ;
  LAYER metal3 ;
  RECT 492.680 646.800 496.220 647.920 ;
  LAYER metal2 ;
  RECT 492.680 646.800 496.220 647.920 ;
  LAYER metal1 ;
  RECT 492.680 646.800 496.220 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 479.040 646.800 482.580 647.920 ;
  LAYER metal4 ;
  RECT 479.040 646.800 482.580 647.920 ;
  LAYER metal3 ;
  RECT 479.040 646.800 482.580 647.920 ;
  LAYER metal2 ;
  RECT 479.040 646.800 482.580 647.920 ;
  LAYER metal1 ;
  RECT 479.040 646.800 482.580 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 465.400 646.800 468.940 647.920 ;
  LAYER metal4 ;
  RECT 465.400 646.800 468.940 647.920 ;
  LAYER metal3 ;
  RECT 465.400 646.800 468.940 647.920 ;
  LAYER metal2 ;
  RECT 465.400 646.800 468.940 647.920 ;
  LAYER metal1 ;
  RECT 465.400 646.800 468.940 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 452.380 646.800 455.920 647.920 ;
  LAYER metal4 ;
  RECT 452.380 646.800 455.920 647.920 ;
  LAYER metal3 ;
  RECT 452.380 646.800 455.920 647.920 ;
  LAYER metal2 ;
  RECT 452.380 646.800 455.920 647.920 ;
  LAYER metal1 ;
  RECT 452.380 646.800 455.920 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 385.420 646.800 388.960 647.920 ;
  LAYER metal4 ;
  RECT 385.420 646.800 388.960 647.920 ;
  LAYER metal3 ;
  RECT 385.420 646.800 388.960 647.920 ;
  LAYER metal2 ;
  RECT 385.420 646.800 388.960 647.920 ;
  LAYER metal1 ;
  RECT 385.420 646.800 388.960 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 376.740 646.800 380.280 647.920 ;
  LAYER metal4 ;
  RECT 376.740 646.800 380.280 647.920 ;
  LAYER metal3 ;
  RECT 376.740 646.800 380.280 647.920 ;
  LAYER metal2 ;
  RECT 376.740 646.800 380.280 647.920 ;
  LAYER metal1 ;
  RECT 376.740 646.800 380.280 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 332.720 646.800 336.260 647.920 ;
  LAYER metal4 ;
  RECT 332.720 646.800 336.260 647.920 ;
  LAYER metal3 ;
  RECT 332.720 646.800 336.260 647.920 ;
  LAYER metal2 ;
  RECT 332.720 646.800 336.260 647.920 ;
  LAYER metal1 ;
  RECT 332.720 646.800 336.260 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 306.680 646.800 310.220 647.920 ;
  LAYER metal4 ;
  RECT 306.680 646.800 310.220 647.920 ;
  LAYER metal3 ;
  RECT 306.680 646.800 310.220 647.920 ;
  LAYER metal2 ;
  RECT 306.680 646.800 310.220 647.920 ;
  LAYER metal1 ;
  RECT 306.680 646.800 310.220 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 298.000 646.800 301.540 647.920 ;
  LAYER metal4 ;
  RECT 298.000 646.800 301.540 647.920 ;
  LAYER metal3 ;
  RECT 298.000 646.800 301.540 647.920 ;
  LAYER metal2 ;
  RECT 298.000 646.800 301.540 647.920 ;
  LAYER metal1 ;
  RECT 298.000 646.800 301.540 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 278.780 646.800 282.320 647.920 ;
  LAYER metal4 ;
  RECT 278.780 646.800 282.320 647.920 ;
  LAYER metal3 ;
  RECT 278.780 646.800 282.320 647.920 ;
  LAYER metal2 ;
  RECT 278.780 646.800 282.320 647.920 ;
  LAYER metal1 ;
  RECT 278.780 646.800 282.320 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 216.780 646.800 220.320 647.920 ;
  LAYER metal4 ;
  RECT 216.780 646.800 220.320 647.920 ;
  LAYER metal3 ;
  RECT 216.780 646.800 220.320 647.920 ;
  LAYER metal2 ;
  RECT 216.780 646.800 220.320 647.920 ;
  LAYER metal1 ;
  RECT 216.780 646.800 220.320 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 203.140 646.800 206.680 647.920 ;
  LAYER metal4 ;
  RECT 203.140 646.800 206.680 647.920 ;
  LAYER metal3 ;
  RECT 203.140 646.800 206.680 647.920 ;
  LAYER metal2 ;
  RECT 203.140 646.800 206.680 647.920 ;
  LAYER metal1 ;
  RECT 203.140 646.800 206.680 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 189.500 646.800 193.040 647.920 ;
  LAYER metal4 ;
  RECT 189.500 646.800 193.040 647.920 ;
  LAYER metal3 ;
  RECT 189.500 646.800 193.040 647.920 ;
  LAYER metal2 ;
  RECT 189.500 646.800 193.040 647.920 ;
  LAYER metal1 ;
  RECT 189.500 646.800 193.040 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 176.480 646.800 180.020 647.920 ;
  LAYER metal4 ;
  RECT 176.480 646.800 180.020 647.920 ;
  LAYER metal3 ;
  RECT 176.480 646.800 180.020 647.920 ;
  LAYER metal2 ;
  RECT 176.480 646.800 180.020 647.920 ;
  LAYER metal1 ;
  RECT 176.480 646.800 180.020 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 162.840 646.800 166.380 647.920 ;
  LAYER metal4 ;
  RECT 162.840 646.800 166.380 647.920 ;
  LAYER metal3 ;
  RECT 162.840 646.800 166.380 647.920 ;
  LAYER metal2 ;
  RECT 162.840 646.800 166.380 647.920 ;
  LAYER metal1 ;
  RECT 162.840 646.800 166.380 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 149.200 646.800 152.740 647.920 ;
  LAYER metal4 ;
  RECT 149.200 646.800 152.740 647.920 ;
  LAYER metal3 ;
  RECT 149.200 646.800 152.740 647.920 ;
  LAYER metal2 ;
  RECT 149.200 646.800 152.740 647.920 ;
  LAYER metal1 ;
  RECT 149.200 646.800 152.740 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 82.240 646.800 85.780 647.920 ;
  LAYER metal4 ;
  RECT 82.240 646.800 85.780 647.920 ;
  LAYER metal3 ;
  RECT 82.240 646.800 85.780 647.920 ;
  LAYER metal2 ;
  RECT 82.240 646.800 85.780 647.920 ;
  LAYER metal1 ;
  RECT 82.240 646.800 85.780 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 68.600 646.800 72.140 647.920 ;
  LAYER metal4 ;
  RECT 68.600 646.800 72.140 647.920 ;
  LAYER metal3 ;
  RECT 68.600 646.800 72.140 647.920 ;
  LAYER metal2 ;
  RECT 68.600 646.800 72.140 647.920 ;
  LAYER metal1 ;
  RECT 68.600 646.800 72.140 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 54.960 646.800 58.500 647.920 ;
  LAYER metal4 ;
  RECT 54.960 646.800 58.500 647.920 ;
  LAYER metal3 ;
  RECT 54.960 646.800 58.500 647.920 ;
  LAYER metal2 ;
  RECT 54.960 646.800 58.500 647.920 ;
  LAYER metal1 ;
  RECT 54.960 646.800 58.500 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 41.940 646.800 45.480 647.920 ;
  LAYER metal4 ;
  RECT 41.940 646.800 45.480 647.920 ;
  LAYER metal3 ;
  RECT 41.940 646.800 45.480 647.920 ;
  LAYER metal2 ;
  RECT 41.940 646.800 45.480 647.920 ;
  LAYER metal1 ;
  RECT 41.940 646.800 45.480 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 28.300 646.800 31.840 647.920 ;
  LAYER metal4 ;
  RECT 28.300 646.800 31.840 647.920 ;
  LAYER metal3 ;
  RECT 28.300 646.800 31.840 647.920 ;
  LAYER metal2 ;
  RECT 28.300 646.800 31.840 647.920 ;
  LAYER metal1 ;
  RECT 28.300 646.800 31.840 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 14.660 646.800 18.200 647.920 ;
  LAYER metal4 ;
  RECT 14.660 646.800 18.200 647.920 ;
  LAYER metal3 ;
  RECT 14.660 646.800 18.200 647.920 ;
  LAYER metal2 ;
  RECT 14.660 646.800 18.200 647.920 ;
  LAYER metal1 ;
  RECT 14.660 646.800 18.200 647.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 653.880 0.000 657.420 1.120 ;
  LAYER metal4 ;
  RECT 653.880 0.000 657.420 1.120 ;
  LAYER metal3 ;
  RECT 653.880 0.000 657.420 1.120 ;
  LAYER metal2 ;
  RECT 653.880 0.000 657.420 1.120 ;
  LAYER metal1 ;
  RECT 653.880 0.000 657.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 640.240 0.000 643.780 1.120 ;
  LAYER metal4 ;
  RECT 640.240 0.000 643.780 1.120 ;
  LAYER metal3 ;
  RECT 640.240 0.000 643.780 1.120 ;
  LAYER metal2 ;
  RECT 640.240 0.000 643.780 1.120 ;
  LAYER metal1 ;
  RECT 640.240 0.000 643.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 627.220 0.000 630.760 1.120 ;
  LAYER metal4 ;
  RECT 627.220 0.000 630.760 1.120 ;
  LAYER metal3 ;
  RECT 627.220 0.000 630.760 1.120 ;
  LAYER metal2 ;
  RECT 627.220 0.000 630.760 1.120 ;
  LAYER metal1 ;
  RECT 627.220 0.000 630.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 613.580 0.000 617.120 1.120 ;
  LAYER metal4 ;
  RECT 613.580 0.000 617.120 1.120 ;
  LAYER metal3 ;
  RECT 613.580 0.000 617.120 1.120 ;
  LAYER metal2 ;
  RECT 613.580 0.000 617.120 1.120 ;
  LAYER metal1 ;
  RECT 613.580 0.000 617.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 599.940 0.000 603.480 1.120 ;
  LAYER metal4 ;
  RECT 599.940 0.000 603.480 1.120 ;
  LAYER metal3 ;
  RECT 599.940 0.000 603.480 1.120 ;
  LAYER metal2 ;
  RECT 599.940 0.000 603.480 1.120 ;
  LAYER metal1 ;
  RECT 599.940 0.000 603.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 586.920 0.000 590.460 1.120 ;
  LAYER metal4 ;
  RECT 586.920 0.000 590.460 1.120 ;
  LAYER metal3 ;
  RECT 586.920 0.000 590.460 1.120 ;
  LAYER metal2 ;
  RECT 586.920 0.000 590.460 1.120 ;
  LAYER metal1 ;
  RECT 586.920 0.000 590.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 519.340 0.000 522.880 1.120 ;
  LAYER metal4 ;
  RECT 519.340 0.000 522.880 1.120 ;
  LAYER metal3 ;
  RECT 519.340 0.000 522.880 1.120 ;
  LAYER metal2 ;
  RECT 519.340 0.000 522.880 1.120 ;
  LAYER metal1 ;
  RECT 519.340 0.000 522.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 506.320 0.000 509.860 1.120 ;
  LAYER metal4 ;
  RECT 506.320 0.000 509.860 1.120 ;
  LAYER metal3 ;
  RECT 506.320 0.000 509.860 1.120 ;
  LAYER metal2 ;
  RECT 506.320 0.000 509.860 1.120 ;
  LAYER metal1 ;
  RECT 506.320 0.000 509.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 492.680 0.000 496.220 1.120 ;
  LAYER metal4 ;
  RECT 492.680 0.000 496.220 1.120 ;
  LAYER metal3 ;
  RECT 492.680 0.000 496.220 1.120 ;
  LAYER metal2 ;
  RECT 492.680 0.000 496.220 1.120 ;
  LAYER metal1 ;
  RECT 492.680 0.000 496.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 479.040 0.000 482.580 1.120 ;
  LAYER metal4 ;
  RECT 479.040 0.000 482.580 1.120 ;
  LAYER metal3 ;
  RECT 479.040 0.000 482.580 1.120 ;
  LAYER metal2 ;
  RECT 479.040 0.000 482.580 1.120 ;
  LAYER metal1 ;
  RECT 479.040 0.000 482.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 465.400 0.000 468.940 1.120 ;
  LAYER metal4 ;
  RECT 465.400 0.000 468.940 1.120 ;
  LAYER metal3 ;
  RECT 465.400 0.000 468.940 1.120 ;
  LAYER metal2 ;
  RECT 465.400 0.000 468.940 1.120 ;
  LAYER metal1 ;
  RECT 465.400 0.000 468.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 452.380 0.000 455.920 1.120 ;
  LAYER metal4 ;
  RECT 452.380 0.000 455.920 1.120 ;
  LAYER metal3 ;
  RECT 452.380 0.000 455.920 1.120 ;
  LAYER metal2 ;
  RECT 452.380 0.000 455.920 1.120 ;
  LAYER metal1 ;
  RECT 452.380 0.000 455.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 385.420 0.000 388.960 1.120 ;
  LAYER metal4 ;
  RECT 385.420 0.000 388.960 1.120 ;
  LAYER metal3 ;
  RECT 385.420 0.000 388.960 1.120 ;
  LAYER metal2 ;
  RECT 385.420 0.000 388.960 1.120 ;
  LAYER metal1 ;
  RECT 385.420 0.000 388.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 376.740 0.000 380.280 1.120 ;
  LAYER metal4 ;
  RECT 376.740 0.000 380.280 1.120 ;
  LAYER metal3 ;
  RECT 376.740 0.000 380.280 1.120 ;
  LAYER metal2 ;
  RECT 376.740 0.000 380.280 1.120 ;
  LAYER metal1 ;
  RECT 376.740 0.000 380.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 332.720 0.000 336.260 1.120 ;
  LAYER metal4 ;
  RECT 332.720 0.000 336.260 1.120 ;
  LAYER metal3 ;
  RECT 332.720 0.000 336.260 1.120 ;
  LAYER metal2 ;
  RECT 332.720 0.000 336.260 1.120 ;
  LAYER metal1 ;
  RECT 332.720 0.000 336.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 306.680 0.000 310.220 1.120 ;
  LAYER metal4 ;
  RECT 306.680 0.000 310.220 1.120 ;
  LAYER metal3 ;
  RECT 306.680 0.000 310.220 1.120 ;
  LAYER metal2 ;
  RECT 306.680 0.000 310.220 1.120 ;
  LAYER metal1 ;
  RECT 306.680 0.000 310.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 298.000 0.000 301.540 1.120 ;
  LAYER metal4 ;
  RECT 298.000 0.000 301.540 1.120 ;
  LAYER metal3 ;
  RECT 298.000 0.000 301.540 1.120 ;
  LAYER metal2 ;
  RECT 298.000 0.000 301.540 1.120 ;
  LAYER metal1 ;
  RECT 298.000 0.000 301.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 278.780 0.000 282.320 1.120 ;
  LAYER metal4 ;
  RECT 278.780 0.000 282.320 1.120 ;
  LAYER metal3 ;
  RECT 278.780 0.000 282.320 1.120 ;
  LAYER metal2 ;
  RECT 278.780 0.000 282.320 1.120 ;
  LAYER metal1 ;
  RECT 278.780 0.000 282.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal4 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal3 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal2 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal1 ;
  RECT 216.780 0.000 220.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal4 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal3 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal2 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal1 ;
  RECT 203.140 0.000 206.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal4 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal3 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal2 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal1 ;
  RECT 189.500 0.000 193.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal4 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal3 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal2 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal1 ;
  RECT 176.480 0.000 180.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal4 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal3 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal2 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal1 ;
  RECT 162.840 0.000 166.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal4 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal3 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal2 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal1 ;
  RECT 149.200 0.000 152.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal4 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal3 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal2 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal1 ;
  RECT 82.240 0.000 85.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal4 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal3 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal2 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal1 ;
  RECT 68.600 0.000 72.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal4 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal3 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal2 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal1 ;
  RECT 54.960 0.000 58.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal4 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal3 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal2 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal1 ;
  RECT 41.940 0.000 45.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal4 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal3 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal2 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal1 ;
  RECT 28.300 0.000 31.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal4 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal3 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal2 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal1 ;
  RECT 14.660 0.000 18.200 1.120 ;
 END
END GND
PIN DIB19
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 651.680 646.800 652.800 647.920 ;
  LAYER metal4 ;
  RECT 651.680 646.800 652.800 647.920 ;
  LAYER metal3 ;
  RECT 651.680 646.800 652.800 647.920 ;
  LAYER metal2 ;
  RECT 651.680 646.800 652.800 647.920 ;
  LAYER metal1 ;
  RECT 651.680 646.800 652.800 647.920 ;
 END
END DIB19
PIN DOB19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 638.040 646.800 639.160 647.920 ;
  LAYER metal4 ;
  RECT 638.040 646.800 639.160 647.920 ;
  LAYER metal3 ;
  RECT 638.040 646.800 639.160 647.920 ;
  LAYER metal2 ;
  RECT 638.040 646.800 639.160 647.920 ;
  LAYER metal1 ;
  RECT 638.040 646.800 639.160 647.920 ;
 END
END DOB19
PIN DIB18
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 625.020 646.800 626.140 647.920 ;
  LAYER metal4 ;
  RECT 625.020 646.800 626.140 647.920 ;
  LAYER metal3 ;
  RECT 625.020 646.800 626.140 647.920 ;
  LAYER metal2 ;
  RECT 625.020 646.800 626.140 647.920 ;
  LAYER metal1 ;
  RECT 625.020 646.800 626.140 647.920 ;
 END
END DIB18
PIN DOB18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 611.380 646.800 612.500 647.920 ;
  LAYER metal4 ;
  RECT 611.380 646.800 612.500 647.920 ;
  LAYER metal3 ;
  RECT 611.380 646.800 612.500 647.920 ;
  LAYER metal2 ;
  RECT 611.380 646.800 612.500 647.920 ;
  LAYER metal1 ;
  RECT 611.380 646.800 612.500 647.920 ;
 END
END DOB18
PIN DIB17
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 597.740 646.800 598.860 647.920 ;
  LAYER metal4 ;
  RECT 597.740 646.800 598.860 647.920 ;
  LAYER metal3 ;
  RECT 597.740 646.800 598.860 647.920 ;
  LAYER metal2 ;
  RECT 597.740 646.800 598.860 647.920 ;
  LAYER metal1 ;
  RECT 597.740 646.800 598.860 647.920 ;
 END
END DIB17
PIN DOB17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 584.720 646.800 585.840 647.920 ;
  LAYER metal4 ;
  RECT 584.720 646.800 585.840 647.920 ;
  LAYER metal3 ;
  RECT 584.720 646.800 585.840 647.920 ;
  LAYER metal2 ;
  RECT 584.720 646.800 585.840 647.920 ;
  LAYER metal1 ;
  RECT 584.720 646.800 585.840 647.920 ;
 END
END DOB17
PIN DIB16
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 571.080 646.800 572.200 647.920 ;
  LAYER metal4 ;
  RECT 571.080 646.800 572.200 647.920 ;
  LAYER metal3 ;
  RECT 571.080 646.800 572.200 647.920 ;
  LAYER metal2 ;
  RECT 571.080 646.800 572.200 647.920 ;
  LAYER metal1 ;
  RECT 571.080 646.800 572.200 647.920 ;
 END
END DIB16
PIN DOB16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 557.440 646.800 558.560 647.920 ;
  LAYER metal4 ;
  RECT 557.440 646.800 558.560 647.920 ;
  LAYER metal3 ;
  RECT 557.440 646.800 558.560 647.920 ;
  LAYER metal2 ;
  RECT 557.440 646.800 558.560 647.920 ;
  LAYER metal1 ;
  RECT 557.440 646.800 558.560 647.920 ;
 END
END DOB16
PIN DIB15
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 544.420 646.800 545.540 647.920 ;
  LAYER metal4 ;
  RECT 544.420 646.800 545.540 647.920 ;
  LAYER metal3 ;
  RECT 544.420 646.800 545.540 647.920 ;
  LAYER metal2 ;
  RECT 544.420 646.800 545.540 647.920 ;
  LAYER metal1 ;
  RECT 544.420 646.800 545.540 647.920 ;
 END
END DIB15
PIN DOB15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 530.780 646.800 531.900 647.920 ;
  LAYER metal4 ;
  RECT 530.780 646.800 531.900 647.920 ;
  LAYER metal3 ;
  RECT 530.780 646.800 531.900 647.920 ;
  LAYER metal2 ;
  RECT 530.780 646.800 531.900 647.920 ;
  LAYER metal1 ;
  RECT 530.780 646.800 531.900 647.920 ;
 END
END DOB15
PIN DIB14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 517.140 646.800 518.260 647.920 ;
  LAYER metal4 ;
  RECT 517.140 646.800 518.260 647.920 ;
  LAYER metal3 ;
  RECT 517.140 646.800 518.260 647.920 ;
  LAYER metal2 ;
  RECT 517.140 646.800 518.260 647.920 ;
  LAYER metal1 ;
  RECT 517.140 646.800 518.260 647.920 ;
 END
END DIB14
PIN DOB14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 504.120 646.800 505.240 647.920 ;
  LAYER metal4 ;
  RECT 504.120 646.800 505.240 647.920 ;
  LAYER metal3 ;
  RECT 504.120 646.800 505.240 647.920 ;
  LAYER metal2 ;
  RECT 504.120 646.800 505.240 647.920 ;
  LAYER metal1 ;
  RECT 504.120 646.800 505.240 647.920 ;
 END
END DOB14
PIN DIB13
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 490.480 646.800 491.600 647.920 ;
  LAYER metal4 ;
  RECT 490.480 646.800 491.600 647.920 ;
  LAYER metal3 ;
  RECT 490.480 646.800 491.600 647.920 ;
  LAYER metal2 ;
  RECT 490.480 646.800 491.600 647.920 ;
  LAYER metal1 ;
  RECT 490.480 646.800 491.600 647.920 ;
 END
END DIB13
PIN DOB13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 476.840 646.800 477.960 647.920 ;
  LAYER metal4 ;
  RECT 476.840 646.800 477.960 647.920 ;
  LAYER metal3 ;
  RECT 476.840 646.800 477.960 647.920 ;
  LAYER metal2 ;
  RECT 476.840 646.800 477.960 647.920 ;
  LAYER metal1 ;
  RECT 476.840 646.800 477.960 647.920 ;
 END
END DOB13
PIN DIB12
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 463.200 646.800 464.320 647.920 ;
  LAYER metal4 ;
  RECT 463.200 646.800 464.320 647.920 ;
  LAYER metal3 ;
  RECT 463.200 646.800 464.320 647.920 ;
  LAYER metal2 ;
  RECT 463.200 646.800 464.320 647.920 ;
  LAYER metal1 ;
  RECT 463.200 646.800 464.320 647.920 ;
 END
END DIB12
PIN DOB12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 450.180 646.800 451.300 647.920 ;
  LAYER metal4 ;
  RECT 450.180 646.800 451.300 647.920 ;
  LAYER metal3 ;
  RECT 450.180 646.800 451.300 647.920 ;
  LAYER metal2 ;
  RECT 450.180 646.800 451.300 647.920 ;
  LAYER metal1 ;
  RECT 450.180 646.800 451.300 647.920 ;
 END
END DOB12
PIN DIB11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 436.540 646.800 437.660 647.920 ;
  LAYER metal4 ;
  RECT 436.540 646.800 437.660 647.920 ;
  LAYER metal3 ;
  RECT 436.540 646.800 437.660 647.920 ;
  LAYER metal2 ;
  RECT 436.540 646.800 437.660 647.920 ;
  LAYER metal1 ;
  RECT 436.540 646.800 437.660 647.920 ;
 END
END DIB11
PIN DOB11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 422.900 646.800 424.020 647.920 ;
  LAYER metal4 ;
  RECT 422.900 646.800 424.020 647.920 ;
  LAYER metal3 ;
  RECT 422.900 646.800 424.020 647.920 ;
  LAYER metal2 ;
  RECT 422.900 646.800 424.020 647.920 ;
  LAYER metal1 ;
  RECT 422.900 646.800 424.020 647.920 ;
 END
END DOB11
PIN DIB10
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 409.880 646.800 411.000 647.920 ;
  LAYER metal4 ;
  RECT 409.880 646.800 411.000 647.920 ;
  LAYER metal3 ;
  RECT 409.880 646.800 411.000 647.920 ;
  LAYER metal2 ;
  RECT 409.880 646.800 411.000 647.920 ;
  LAYER metal1 ;
  RECT 409.880 646.800 411.000 647.920 ;
 END
END DIB10
PIN DOB10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 396.240 646.800 397.360 647.920 ;
  LAYER metal4 ;
  RECT 396.240 646.800 397.360 647.920 ;
  LAYER metal3 ;
  RECT 396.240 646.800 397.360 647.920 ;
  LAYER metal2 ;
  RECT 396.240 646.800 397.360 647.920 ;
  LAYER metal1 ;
  RECT 396.240 646.800 397.360 647.920 ;
 END
END DOB10
PIN CKB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 374.540 646.800 375.660 647.920 ;
  LAYER metal4 ;
  RECT 374.540 646.800 375.660 647.920 ;
  LAYER metal3 ;
  RECT 374.540 646.800 375.660 647.920 ;
  LAYER metal2 ;
  RECT 374.540 646.800 375.660 647.920 ;
  LAYER metal1 ;
  RECT 374.540 646.800 375.660 647.920 ;
 END
END CKB
PIN CSB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 372.060 646.800 373.180 647.920 ;
  LAYER metal4 ;
  RECT 372.060 646.800 373.180 647.920 ;
  LAYER metal3 ;
  RECT 372.060 646.800 373.180 647.920 ;
  LAYER metal2 ;
  RECT 372.060 646.800 373.180 647.920 ;
  LAYER metal1 ;
  RECT 372.060 646.800 373.180 647.920 ;
 END
END CSB
PIN WEBN
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 370.200 646.800 371.320 647.920 ;
  LAYER metal4 ;
  RECT 370.200 646.800 371.320 647.920 ;
  LAYER metal3 ;
  RECT 370.200 646.800 371.320 647.920 ;
  LAYER metal2 ;
  RECT 370.200 646.800 371.320 647.920 ;
  LAYER metal1 ;
  RECT 370.200 646.800 371.320 647.920 ;
 END
END WEBN
PIN B2
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 366.480 646.800 367.600 647.920 ;
  LAYER metal4 ;
  RECT 366.480 646.800 367.600 647.920 ;
  LAYER metal3 ;
  RECT 366.480 646.800 367.600 647.920 ;
  LAYER metal2 ;
  RECT 366.480 646.800 367.600 647.920 ;
  LAYER metal1 ;
  RECT 366.480 646.800 367.600 647.920 ;
 END
END B2
PIN OEB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 362.760 646.800 363.880 647.920 ;
  LAYER metal4 ;
  RECT 362.760 646.800 363.880 647.920 ;
  LAYER metal3 ;
  RECT 362.760 646.800 363.880 647.920 ;
  LAYER metal2 ;
  RECT 362.760 646.800 363.880 647.920 ;
  LAYER metal1 ;
  RECT 362.760 646.800 363.880 647.920 ;
 END
END OEB
PIN B1
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 360.900 646.800 362.020 647.920 ;
  LAYER metal4 ;
  RECT 360.900 646.800 362.020 647.920 ;
  LAYER metal3 ;
  RECT 360.900 646.800 362.020 647.920 ;
  LAYER metal2 ;
  RECT 360.900 646.800 362.020 647.920 ;
  LAYER metal1 ;
  RECT 360.900 646.800 362.020 647.920 ;
 END
END B1
PIN B0
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 359.040 646.800 360.160 647.920 ;
  LAYER metal4 ;
  RECT 359.040 646.800 360.160 647.920 ;
  LAYER metal3 ;
  RECT 359.040 646.800 360.160 647.920 ;
  LAYER metal2 ;
  RECT 359.040 646.800 360.160 647.920 ;
  LAYER metal1 ;
  RECT 359.040 646.800 360.160 647.920 ;
 END
END B0
PIN B5
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 350.360 646.800 351.480 647.920 ;
  LAYER metal4 ;
  RECT 350.360 646.800 351.480 647.920 ;
  LAYER metal3 ;
  RECT 350.360 646.800 351.480 647.920 ;
  LAYER metal2 ;
  RECT 350.360 646.800 351.480 647.920 ;
  LAYER metal1 ;
  RECT 350.360 646.800 351.480 647.920 ;
 END
END B5
PIN B4
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 344.780 646.800 345.900 647.920 ;
  LAYER metal4 ;
  RECT 344.780 646.800 345.900 647.920 ;
  LAYER metal3 ;
  RECT 344.780 646.800 345.900 647.920 ;
  LAYER metal2 ;
  RECT 344.780 646.800 345.900 647.920 ;
  LAYER metal1 ;
  RECT 344.780 646.800 345.900 647.920 ;
 END
END B4
PIN B3
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 339.200 646.800 340.320 647.920 ;
  LAYER metal4 ;
  RECT 339.200 646.800 340.320 647.920 ;
  LAYER metal3 ;
  RECT 339.200 646.800 340.320 647.920 ;
  LAYER metal2 ;
  RECT 339.200 646.800 340.320 647.920 ;
  LAYER metal1 ;
  RECT 339.200 646.800 340.320 647.920 ;
 END
END B3
PIN B8
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 326.180 646.800 327.300 647.920 ;
  LAYER metal4 ;
  RECT 326.180 646.800 327.300 647.920 ;
  LAYER metal3 ;
  RECT 326.180 646.800 327.300 647.920 ;
  LAYER metal2 ;
  RECT 326.180 646.800 327.300 647.920 ;
  LAYER metal1 ;
  RECT 326.180 646.800 327.300 647.920 ;
 END
END B8
PIN B7
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 320.600 646.800 321.720 647.920 ;
  LAYER metal4 ;
  RECT 320.600 646.800 321.720 647.920 ;
  LAYER metal3 ;
  RECT 320.600 646.800 321.720 647.920 ;
  LAYER metal2 ;
  RECT 320.600 646.800 321.720 647.920 ;
  LAYER metal1 ;
  RECT 320.600 646.800 321.720 647.920 ;
 END
END B7
PIN B6
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 314.400 646.800 315.520 647.920 ;
  LAYER metal4 ;
  RECT 314.400 646.800 315.520 647.920 ;
  LAYER metal3 ;
  RECT 314.400 646.800 315.520 647.920 ;
  LAYER metal2 ;
  RECT 314.400 646.800 315.520 647.920 ;
  LAYER metal1 ;
  RECT 314.400 646.800 315.520 647.920 ;
 END
END B6
PIN B10
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 295.800 646.800 296.920 647.920 ;
  LAYER metal4 ;
  RECT 295.800 646.800 296.920 647.920 ;
  LAYER metal3 ;
  RECT 295.800 646.800 296.920 647.920 ;
  LAYER metal2 ;
  RECT 295.800 646.800 296.920 647.920 ;
  LAYER metal1 ;
  RECT 295.800 646.800 296.920 647.920 ;
 END
END B10
PIN B9
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 290.220 646.800 291.340 647.920 ;
  LAYER metal4 ;
  RECT 290.220 646.800 291.340 647.920 ;
  LAYER metal3 ;
  RECT 290.220 646.800 291.340 647.920 ;
  LAYER metal2 ;
  RECT 290.220 646.800 291.340 647.920 ;
  LAYER metal1 ;
  RECT 290.220 646.800 291.340 647.920 ;
 END
END B9
PIN DIB9
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 267.900 646.800 269.020 647.920 ;
  LAYER metal4 ;
  RECT 267.900 646.800 269.020 647.920 ;
  LAYER metal3 ;
  RECT 267.900 646.800 269.020 647.920 ;
  LAYER metal2 ;
  RECT 267.900 646.800 269.020 647.920 ;
  LAYER metal1 ;
  RECT 267.900 646.800 269.020 647.920 ;
 END
END DIB9
PIN DOB9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 254.880 646.800 256.000 647.920 ;
  LAYER metal4 ;
  RECT 254.880 646.800 256.000 647.920 ;
  LAYER metal3 ;
  RECT 254.880 646.800 256.000 647.920 ;
  LAYER metal2 ;
  RECT 254.880 646.800 256.000 647.920 ;
  LAYER metal1 ;
  RECT 254.880 646.800 256.000 647.920 ;
 END
END DOB9
PIN DIB8
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 241.240 646.800 242.360 647.920 ;
  LAYER metal4 ;
  RECT 241.240 646.800 242.360 647.920 ;
  LAYER metal3 ;
  RECT 241.240 646.800 242.360 647.920 ;
  LAYER metal2 ;
  RECT 241.240 646.800 242.360 647.920 ;
  LAYER metal1 ;
  RECT 241.240 646.800 242.360 647.920 ;
 END
END DIB8
PIN DOB8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 227.600 646.800 228.720 647.920 ;
  LAYER metal4 ;
  RECT 227.600 646.800 228.720 647.920 ;
  LAYER metal3 ;
  RECT 227.600 646.800 228.720 647.920 ;
  LAYER metal2 ;
  RECT 227.600 646.800 228.720 647.920 ;
  LAYER metal1 ;
  RECT 227.600 646.800 228.720 647.920 ;
 END
END DOB8
PIN DIB7
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 214.580 646.800 215.700 647.920 ;
  LAYER metal4 ;
  RECT 214.580 646.800 215.700 647.920 ;
  LAYER metal3 ;
  RECT 214.580 646.800 215.700 647.920 ;
  LAYER metal2 ;
  RECT 214.580 646.800 215.700 647.920 ;
  LAYER metal1 ;
  RECT 214.580 646.800 215.700 647.920 ;
 END
END DIB7
PIN DOB7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 200.940 646.800 202.060 647.920 ;
  LAYER metal4 ;
  RECT 200.940 646.800 202.060 647.920 ;
  LAYER metal3 ;
  RECT 200.940 646.800 202.060 647.920 ;
  LAYER metal2 ;
  RECT 200.940 646.800 202.060 647.920 ;
  LAYER metal1 ;
  RECT 200.940 646.800 202.060 647.920 ;
 END
END DOB7
PIN DIB6
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 187.300 646.800 188.420 647.920 ;
  LAYER metal4 ;
  RECT 187.300 646.800 188.420 647.920 ;
  LAYER metal3 ;
  RECT 187.300 646.800 188.420 647.920 ;
  LAYER metal2 ;
  RECT 187.300 646.800 188.420 647.920 ;
  LAYER metal1 ;
  RECT 187.300 646.800 188.420 647.920 ;
 END
END DIB6
PIN DOB6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 174.280 646.800 175.400 647.920 ;
  LAYER metal4 ;
  RECT 174.280 646.800 175.400 647.920 ;
  LAYER metal3 ;
  RECT 174.280 646.800 175.400 647.920 ;
  LAYER metal2 ;
  RECT 174.280 646.800 175.400 647.920 ;
  LAYER metal1 ;
  RECT 174.280 646.800 175.400 647.920 ;
 END
END DOB6
PIN DIB5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 160.640 646.800 161.760 647.920 ;
  LAYER metal4 ;
  RECT 160.640 646.800 161.760 647.920 ;
  LAYER metal3 ;
  RECT 160.640 646.800 161.760 647.920 ;
  LAYER metal2 ;
  RECT 160.640 646.800 161.760 647.920 ;
  LAYER metal1 ;
  RECT 160.640 646.800 161.760 647.920 ;
 END
END DIB5
PIN DOB5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 147.000 646.800 148.120 647.920 ;
  LAYER metal4 ;
  RECT 147.000 646.800 148.120 647.920 ;
  LAYER metal3 ;
  RECT 147.000 646.800 148.120 647.920 ;
  LAYER metal2 ;
  RECT 147.000 646.800 148.120 647.920 ;
  LAYER metal1 ;
  RECT 147.000 646.800 148.120 647.920 ;
 END
END DOB5
PIN DIB4
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 133.980 646.800 135.100 647.920 ;
  LAYER metal4 ;
  RECT 133.980 646.800 135.100 647.920 ;
  LAYER metal3 ;
  RECT 133.980 646.800 135.100 647.920 ;
  LAYER metal2 ;
  RECT 133.980 646.800 135.100 647.920 ;
  LAYER metal1 ;
  RECT 133.980 646.800 135.100 647.920 ;
 END
END DIB4
PIN DOB4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 120.340 646.800 121.460 647.920 ;
  LAYER metal4 ;
  RECT 120.340 646.800 121.460 647.920 ;
  LAYER metal3 ;
  RECT 120.340 646.800 121.460 647.920 ;
  LAYER metal2 ;
  RECT 120.340 646.800 121.460 647.920 ;
  LAYER metal1 ;
  RECT 120.340 646.800 121.460 647.920 ;
 END
END DOB4
PIN DIB3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 106.700 646.800 107.820 647.920 ;
  LAYER metal4 ;
  RECT 106.700 646.800 107.820 647.920 ;
  LAYER metal3 ;
  RECT 106.700 646.800 107.820 647.920 ;
  LAYER metal2 ;
  RECT 106.700 646.800 107.820 647.920 ;
  LAYER metal1 ;
  RECT 106.700 646.800 107.820 647.920 ;
 END
END DIB3
PIN DOB3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 93.680 646.800 94.800 647.920 ;
  LAYER metal4 ;
  RECT 93.680 646.800 94.800 647.920 ;
  LAYER metal3 ;
  RECT 93.680 646.800 94.800 647.920 ;
  LAYER metal2 ;
  RECT 93.680 646.800 94.800 647.920 ;
  LAYER metal1 ;
  RECT 93.680 646.800 94.800 647.920 ;
 END
END DOB3
PIN DIB2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 80.040 646.800 81.160 647.920 ;
  LAYER metal4 ;
  RECT 80.040 646.800 81.160 647.920 ;
  LAYER metal3 ;
  RECT 80.040 646.800 81.160 647.920 ;
  LAYER metal2 ;
  RECT 80.040 646.800 81.160 647.920 ;
  LAYER metal1 ;
  RECT 80.040 646.800 81.160 647.920 ;
 END
END DIB2
PIN DOB2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 66.400 646.800 67.520 647.920 ;
  LAYER metal4 ;
  RECT 66.400 646.800 67.520 647.920 ;
  LAYER metal3 ;
  RECT 66.400 646.800 67.520 647.920 ;
  LAYER metal2 ;
  RECT 66.400 646.800 67.520 647.920 ;
  LAYER metal1 ;
  RECT 66.400 646.800 67.520 647.920 ;
 END
END DOB2
PIN DIB1
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 52.760 646.800 53.880 647.920 ;
  LAYER metal4 ;
  RECT 52.760 646.800 53.880 647.920 ;
  LAYER metal3 ;
  RECT 52.760 646.800 53.880 647.920 ;
  LAYER metal2 ;
  RECT 52.760 646.800 53.880 647.920 ;
  LAYER metal1 ;
  RECT 52.760 646.800 53.880 647.920 ;
 END
END DIB1
PIN DOB1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 39.740 646.800 40.860 647.920 ;
  LAYER metal4 ;
  RECT 39.740 646.800 40.860 647.920 ;
  LAYER metal3 ;
  RECT 39.740 646.800 40.860 647.920 ;
  LAYER metal2 ;
  RECT 39.740 646.800 40.860 647.920 ;
  LAYER metal1 ;
  RECT 39.740 646.800 40.860 647.920 ;
 END
END DOB1
PIN DIB0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 26.100 646.800 27.220 647.920 ;
  LAYER metal4 ;
  RECT 26.100 646.800 27.220 647.920 ;
  LAYER metal3 ;
  RECT 26.100 646.800 27.220 647.920 ;
  LAYER metal2 ;
  RECT 26.100 646.800 27.220 647.920 ;
  LAYER metal1 ;
  RECT 26.100 646.800 27.220 647.920 ;
 END
END DIB0
PIN DOB0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 12.460 646.800 13.580 647.920 ;
  LAYER metal4 ;
  RECT 12.460 646.800 13.580 647.920 ;
  LAYER metal3 ;
  RECT 12.460 646.800 13.580 647.920 ;
  LAYER metal2 ;
  RECT 12.460 646.800 13.580 647.920 ;
  LAYER metal1 ;
  RECT 12.460 646.800 13.580 647.920 ;
 END
END DOB0
PIN DIA19
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 651.680 0.000 652.800 1.120 ;
  LAYER metal4 ;
  RECT 651.680 0.000 652.800 1.120 ;
  LAYER metal3 ;
  RECT 651.680 0.000 652.800 1.120 ;
  LAYER metal2 ;
  RECT 651.680 0.000 652.800 1.120 ;
  LAYER metal1 ;
  RECT 651.680 0.000 652.800 1.120 ;
 END
END DIA19
PIN DOA19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 638.040 0.000 639.160 1.120 ;
  LAYER metal4 ;
  RECT 638.040 0.000 639.160 1.120 ;
  LAYER metal3 ;
  RECT 638.040 0.000 639.160 1.120 ;
  LAYER metal2 ;
  RECT 638.040 0.000 639.160 1.120 ;
  LAYER metal1 ;
  RECT 638.040 0.000 639.160 1.120 ;
 END
END DOA19
PIN DIA18
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 625.020 0.000 626.140 1.120 ;
  LAYER metal4 ;
  RECT 625.020 0.000 626.140 1.120 ;
  LAYER metal3 ;
  RECT 625.020 0.000 626.140 1.120 ;
  LAYER metal2 ;
  RECT 625.020 0.000 626.140 1.120 ;
  LAYER metal1 ;
  RECT 625.020 0.000 626.140 1.120 ;
 END
END DIA18
PIN DOA18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 611.380 0.000 612.500 1.120 ;
  LAYER metal4 ;
  RECT 611.380 0.000 612.500 1.120 ;
  LAYER metal3 ;
  RECT 611.380 0.000 612.500 1.120 ;
  LAYER metal2 ;
  RECT 611.380 0.000 612.500 1.120 ;
  LAYER metal1 ;
  RECT 611.380 0.000 612.500 1.120 ;
 END
END DOA18
PIN DIA17
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 597.740 0.000 598.860 1.120 ;
  LAYER metal4 ;
  RECT 597.740 0.000 598.860 1.120 ;
  LAYER metal3 ;
  RECT 597.740 0.000 598.860 1.120 ;
  LAYER metal2 ;
  RECT 597.740 0.000 598.860 1.120 ;
  LAYER metal1 ;
  RECT 597.740 0.000 598.860 1.120 ;
 END
END DIA17
PIN DOA17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 584.720 0.000 585.840 1.120 ;
  LAYER metal4 ;
  RECT 584.720 0.000 585.840 1.120 ;
  LAYER metal3 ;
  RECT 584.720 0.000 585.840 1.120 ;
  LAYER metal2 ;
  RECT 584.720 0.000 585.840 1.120 ;
  LAYER metal1 ;
  RECT 584.720 0.000 585.840 1.120 ;
 END
END DOA17
PIN DIA16
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 571.080 0.000 572.200 1.120 ;
  LAYER metal4 ;
  RECT 571.080 0.000 572.200 1.120 ;
  LAYER metal3 ;
  RECT 571.080 0.000 572.200 1.120 ;
  LAYER metal2 ;
  RECT 571.080 0.000 572.200 1.120 ;
  LAYER metal1 ;
  RECT 571.080 0.000 572.200 1.120 ;
 END
END DIA16
PIN DOA16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 557.440 0.000 558.560 1.120 ;
  LAYER metal4 ;
  RECT 557.440 0.000 558.560 1.120 ;
  LAYER metal3 ;
  RECT 557.440 0.000 558.560 1.120 ;
  LAYER metal2 ;
  RECT 557.440 0.000 558.560 1.120 ;
  LAYER metal1 ;
  RECT 557.440 0.000 558.560 1.120 ;
 END
END DOA16
PIN DIA15
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 544.420 0.000 545.540 1.120 ;
  LAYER metal4 ;
  RECT 544.420 0.000 545.540 1.120 ;
  LAYER metal3 ;
  RECT 544.420 0.000 545.540 1.120 ;
  LAYER metal2 ;
  RECT 544.420 0.000 545.540 1.120 ;
  LAYER metal1 ;
  RECT 544.420 0.000 545.540 1.120 ;
 END
END DIA15
PIN DOA15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER metal4 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER metal3 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER metal2 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER metal1 ;
  RECT 530.780 0.000 531.900 1.120 ;
 END
END DOA15
PIN DIA14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 517.140 0.000 518.260 1.120 ;
  LAYER metal4 ;
  RECT 517.140 0.000 518.260 1.120 ;
  LAYER metal3 ;
  RECT 517.140 0.000 518.260 1.120 ;
  LAYER metal2 ;
  RECT 517.140 0.000 518.260 1.120 ;
  LAYER metal1 ;
  RECT 517.140 0.000 518.260 1.120 ;
 END
END DIA14
PIN DOA14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 504.120 0.000 505.240 1.120 ;
  LAYER metal4 ;
  RECT 504.120 0.000 505.240 1.120 ;
  LAYER metal3 ;
  RECT 504.120 0.000 505.240 1.120 ;
  LAYER metal2 ;
  RECT 504.120 0.000 505.240 1.120 ;
  LAYER metal1 ;
  RECT 504.120 0.000 505.240 1.120 ;
 END
END DOA14
PIN DIA13
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 490.480 0.000 491.600 1.120 ;
  LAYER metal4 ;
  RECT 490.480 0.000 491.600 1.120 ;
  LAYER metal3 ;
  RECT 490.480 0.000 491.600 1.120 ;
  LAYER metal2 ;
  RECT 490.480 0.000 491.600 1.120 ;
  LAYER metal1 ;
  RECT 490.480 0.000 491.600 1.120 ;
 END
END DIA13
PIN DOA13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 476.840 0.000 477.960 1.120 ;
  LAYER metal4 ;
  RECT 476.840 0.000 477.960 1.120 ;
  LAYER metal3 ;
  RECT 476.840 0.000 477.960 1.120 ;
  LAYER metal2 ;
  RECT 476.840 0.000 477.960 1.120 ;
  LAYER metal1 ;
  RECT 476.840 0.000 477.960 1.120 ;
 END
END DOA13
PIN DIA12
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 463.200 0.000 464.320 1.120 ;
  LAYER metal4 ;
  RECT 463.200 0.000 464.320 1.120 ;
  LAYER metal3 ;
  RECT 463.200 0.000 464.320 1.120 ;
  LAYER metal2 ;
  RECT 463.200 0.000 464.320 1.120 ;
  LAYER metal1 ;
  RECT 463.200 0.000 464.320 1.120 ;
 END
END DIA12
PIN DOA12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 450.180 0.000 451.300 1.120 ;
  LAYER metal4 ;
  RECT 450.180 0.000 451.300 1.120 ;
  LAYER metal3 ;
  RECT 450.180 0.000 451.300 1.120 ;
  LAYER metal2 ;
  RECT 450.180 0.000 451.300 1.120 ;
  LAYER metal1 ;
  RECT 450.180 0.000 451.300 1.120 ;
 END
END DOA12
PIN DIA11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 436.540 0.000 437.660 1.120 ;
  LAYER metal4 ;
  RECT 436.540 0.000 437.660 1.120 ;
  LAYER metal3 ;
  RECT 436.540 0.000 437.660 1.120 ;
  LAYER metal2 ;
  RECT 436.540 0.000 437.660 1.120 ;
  LAYER metal1 ;
  RECT 436.540 0.000 437.660 1.120 ;
 END
END DIA11
PIN DOA11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 422.900 0.000 424.020 1.120 ;
  LAYER metal4 ;
  RECT 422.900 0.000 424.020 1.120 ;
  LAYER metal3 ;
  RECT 422.900 0.000 424.020 1.120 ;
  LAYER metal2 ;
  RECT 422.900 0.000 424.020 1.120 ;
  LAYER metal1 ;
  RECT 422.900 0.000 424.020 1.120 ;
 END
END DOA11
PIN DIA10
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 409.880 0.000 411.000 1.120 ;
  LAYER metal4 ;
  RECT 409.880 0.000 411.000 1.120 ;
  LAYER metal3 ;
  RECT 409.880 0.000 411.000 1.120 ;
  LAYER metal2 ;
  RECT 409.880 0.000 411.000 1.120 ;
  LAYER metal1 ;
  RECT 409.880 0.000 411.000 1.120 ;
 END
END DIA10
PIN DOA10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 396.240 0.000 397.360 1.120 ;
  LAYER metal4 ;
  RECT 396.240 0.000 397.360 1.120 ;
  LAYER metal3 ;
  RECT 396.240 0.000 397.360 1.120 ;
  LAYER metal2 ;
  RECT 396.240 0.000 397.360 1.120 ;
  LAYER metal1 ;
  RECT 396.240 0.000 397.360 1.120 ;
 END
END DOA10
PIN CKA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 374.540 0.000 375.660 1.120 ;
  LAYER metal4 ;
  RECT 374.540 0.000 375.660 1.120 ;
  LAYER metal3 ;
  RECT 374.540 0.000 375.660 1.120 ;
  LAYER metal2 ;
  RECT 374.540 0.000 375.660 1.120 ;
  LAYER metal1 ;
  RECT 374.540 0.000 375.660 1.120 ;
 END
END CKA
PIN CSA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 372.060 0.000 373.180 1.120 ;
  LAYER metal4 ;
  RECT 372.060 0.000 373.180 1.120 ;
  LAYER metal3 ;
  RECT 372.060 0.000 373.180 1.120 ;
  LAYER metal2 ;
  RECT 372.060 0.000 373.180 1.120 ;
  LAYER metal1 ;
  RECT 372.060 0.000 373.180 1.120 ;
 END
END CSA
PIN WEAN
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 370.200 0.000 371.320 1.120 ;
  LAYER metal4 ;
  RECT 370.200 0.000 371.320 1.120 ;
  LAYER metal3 ;
  RECT 370.200 0.000 371.320 1.120 ;
  LAYER metal2 ;
  RECT 370.200 0.000 371.320 1.120 ;
  LAYER metal1 ;
  RECT 370.200 0.000 371.320 1.120 ;
 END
END WEAN
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 366.480 0.000 367.600 1.120 ;
  LAYER metal4 ;
  RECT 366.480 0.000 367.600 1.120 ;
  LAYER metal3 ;
  RECT 366.480 0.000 367.600 1.120 ;
  LAYER metal2 ;
  RECT 366.480 0.000 367.600 1.120 ;
  LAYER metal1 ;
  RECT 366.480 0.000 367.600 1.120 ;
 END
END A2
PIN OEA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 362.760 0.000 363.880 1.120 ;
  LAYER metal4 ;
  RECT 362.760 0.000 363.880 1.120 ;
  LAYER metal3 ;
  RECT 362.760 0.000 363.880 1.120 ;
  LAYER metal2 ;
  RECT 362.760 0.000 363.880 1.120 ;
  LAYER metal1 ;
  RECT 362.760 0.000 363.880 1.120 ;
 END
END OEA
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 360.900 0.000 362.020 1.120 ;
  LAYER metal4 ;
  RECT 360.900 0.000 362.020 1.120 ;
  LAYER metal3 ;
  RECT 360.900 0.000 362.020 1.120 ;
  LAYER metal2 ;
  RECT 360.900 0.000 362.020 1.120 ;
  LAYER metal1 ;
  RECT 360.900 0.000 362.020 1.120 ;
 END
END A1
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal4 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal3 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal2 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal1 ;
  RECT 359.040 0.000 360.160 1.120 ;
 END
END A0
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 350.360 0.000 351.480 1.120 ;
  LAYER metal4 ;
  RECT 350.360 0.000 351.480 1.120 ;
  LAYER metal3 ;
  RECT 350.360 0.000 351.480 1.120 ;
  LAYER metal2 ;
  RECT 350.360 0.000 351.480 1.120 ;
  LAYER metal1 ;
  RECT 350.360 0.000 351.480 1.120 ;
 END
END A5
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 344.780 0.000 345.900 1.120 ;
  LAYER metal4 ;
  RECT 344.780 0.000 345.900 1.120 ;
  LAYER metal3 ;
  RECT 344.780 0.000 345.900 1.120 ;
  LAYER metal2 ;
  RECT 344.780 0.000 345.900 1.120 ;
  LAYER metal1 ;
  RECT 344.780 0.000 345.900 1.120 ;
 END
END A4
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 339.200 0.000 340.320 1.120 ;
  LAYER metal4 ;
  RECT 339.200 0.000 340.320 1.120 ;
  LAYER metal3 ;
  RECT 339.200 0.000 340.320 1.120 ;
  LAYER metal2 ;
  RECT 339.200 0.000 340.320 1.120 ;
  LAYER metal1 ;
  RECT 339.200 0.000 340.320 1.120 ;
 END
END A3
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 326.180 0.000 327.300 1.120 ;
  LAYER metal4 ;
  RECT 326.180 0.000 327.300 1.120 ;
  LAYER metal3 ;
  RECT 326.180 0.000 327.300 1.120 ;
  LAYER metal2 ;
  RECT 326.180 0.000 327.300 1.120 ;
  LAYER metal1 ;
  RECT 326.180 0.000 327.300 1.120 ;
 END
END A8
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 320.600 0.000 321.720 1.120 ;
  LAYER metal4 ;
  RECT 320.600 0.000 321.720 1.120 ;
  LAYER metal3 ;
  RECT 320.600 0.000 321.720 1.120 ;
  LAYER metal2 ;
  RECT 320.600 0.000 321.720 1.120 ;
  LAYER metal1 ;
  RECT 320.600 0.000 321.720 1.120 ;
 END
END A7
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 314.400 0.000 315.520 1.120 ;
  LAYER metal4 ;
  RECT 314.400 0.000 315.520 1.120 ;
  LAYER metal3 ;
  RECT 314.400 0.000 315.520 1.120 ;
  LAYER metal2 ;
  RECT 314.400 0.000 315.520 1.120 ;
  LAYER metal1 ;
  RECT 314.400 0.000 315.520 1.120 ;
 END
END A6
PIN A10
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 295.800 0.000 296.920 1.120 ;
  LAYER metal4 ;
  RECT 295.800 0.000 296.920 1.120 ;
  LAYER metal3 ;
  RECT 295.800 0.000 296.920 1.120 ;
  LAYER metal2 ;
  RECT 295.800 0.000 296.920 1.120 ;
  LAYER metal1 ;
  RECT 295.800 0.000 296.920 1.120 ;
 END
END A10
PIN A9
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 290.220 0.000 291.340 1.120 ;
  LAYER metal4 ;
  RECT 290.220 0.000 291.340 1.120 ;
  LAYER metal3 ;
  RECT 290.220 0.000 291.340 1.120 ;
  LAYER metal2 ;
  RECT 290.220 0.000 291.340 1.120 ;
  LAYER metal1 ;
  RECT 290.220 0.000 291.340 1.120 ;
 END
END A9
PIN DIA9
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal4 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal3 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal2 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal1 ;
  RECT 267.900 0.000 269.020 1.120 ;
 END
END DIA9
PIN DOA9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal4 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal3 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal2 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal1 ;
  RECT 254.880 0.000 256.000 1.120 ;
 END
END DOA9
PIN DIA8
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal4 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal3 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal2 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal1 ;
  RECT 241.240 0.000 242.360 1.120 ;
 END
END DIA8
PIN DOA8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal4 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal3 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal2 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal1 ;
  RECT 227.600 0.000 228.720 1.120 ;
 END
END DOA8
PIN DIA7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal4 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal3 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal2 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal1 ;
  RECT 214.580 0.000 215.700 1.120 ;
 END
END DIA7
PIN DOA7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal4 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal3 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal2 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal1 ;
  RECT 200.940 0.000 202.060 1.120 ;
 END
END DOA7
PIN DIA6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal4 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal3 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal2 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal1 ;
  RECT 187.300 0.000 188.420 1.120 ;
 END
END DIA6
PIN DOA6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal4 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal3 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal2 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal1 ;
  RECT 174.280 0.000 175.400 1.120 ;
 END
END DOA6
PIN DIA5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal4 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal3 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal2 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal1 ;
  RECT 160.640 0.000 161.760 1.120 ;
 END
END DIA5
PIN DOA5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal4 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal3 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal2 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal1 ;
  RECT 147.000 0.000 148.120 1.120 ;
 END
END DOA5
PIN DIA4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal4 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal3 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal2 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal1 ;
  RECT 133.980 0.000 135.100 1.120 ;
 END
END DIA4
PIN DOA4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal4 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal3 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal2 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal1 ;
  RECT 120.340 0.000 121.460 1.120 ;
 END
END DOA4
PIN DIA3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DIA3
PIN DOA3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal4 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal3 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal2 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal1 ;
  RECT 93.680 0.000 94.800 1.120 ;
 END
END DOA3
PIN DIA2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal4 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal3 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal2 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal1 ;
  RECT 80.040 0.000 81.160 1.120 ;
 END
END DIA2
PIN DOA2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal4 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal3 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal2 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal1 ;
  RECT 66.400 0.000 67.520 1.120 ;
 END
END DOA2
PIN DIA1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal4 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal3 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal2 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal1 ;
  RECT 52.760 0.000 53.880 1.120 ;
 END
END DIA1
PIN DOA1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal4 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal3 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal2 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal1 ;
  RECT 39.740 0.000 40.860 1.120 ;
 END
END DOA1
PIN DIA0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal4 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal3 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal2 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal1 ;
  RECT 26.100 0.000 27.220 1.120 ;
 END
END DIA0
PIN DOA0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal4 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal3 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal2 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal1 ;
  RECT 12.460 0.000 13.580 1.120 ;
 END
END DOA0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 674.560 647.780 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 674.560 647.780 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 674.560 647.780 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 674.560 647.780 ;
  LAYER via ;
  RECT 0.000 0.140 674.560 647.780 ;
  LAYER via2 ;
  RECT 0.000 0.140 674.560 647.780 ;
  LAYER via3 ;
  RECT 0.000 0.140 674.560 647.780 ;
END
END SRAM_1296X20
END LIBRARY



